`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 2017/12/31 21:04:21
// Design Name: 
// Module Name: color_rom2
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module color_rom2(input ena,input [14:0]addr,output reg [11:0]color);
always@(ena)
begin
if(ena)
begin
color<=12'bz;
end
else
begin
case(addr)
15'b0000100111010100011 : color = 12'he73;
15'b0000100111010100100 : color = 12'he73;
15'b0000100111010100101 : color = 12'he73;
15'b0000100111010100110 : color = 12'he73;
15'b0000100111010100111 : color = 12'he73;
15'b0000100111010101000 : color = 12'he73;
15'b0000100111010101001 : color = 12'he73;
15'b0000100111010101010 : color = 12'he73;
15'b0000100111010101011 : color = 12'he73;
15'b0000100111010101100 : color = 12'he73;
15'b0000100111010101101 : color = 12'he73;
15'b0000100111010101110 : color = 12'he73;
15'b0000100111010101111 : color = 12'he73;
15'b0000100111010110000 : color = 12'he73;
15'b0000100111010110001 : color = 12'he73;
15'b0000100111010110010 : color = 12'he73;
15'b0000100111010110011 : color = 12'he73;
15'b0000100111010110100 : color = 12'he73;
15'b0000100111010110101 : color = 12'he73;
15'b0000100111010110110 : color = 12'he73;
15'b0000100111010110111 : color = 12'he73;
15'b0000100111010111000 : color = 12'he73;
15'b0000100111010111001 : color = 12'he73;
15'b0000100111010111010 : color = 12'he73;
15'b0000100111010111011 : color = 12'he73;
15'b0000100111010111100 : color = 12'he73;
15'b0000100111010111101 : color = 12'he73;
15'b0000100111010111110 : color = 12'he73;
15'b0000100111010111111 : color = 12'he73;
15'b0000100111011000000 : color = 12'he73;
15'b0000100111011000001 : color = 12'he73;
15'b0000100111011000010 : color = 12'he73;
15'b0000100111011000011 : color = 12'he73;
15'b0000100111011000100 : color = 12'he73;
15'b0000100111011000101 : color = 12'he73;
15'b0000100111011000110 : color = 12'he73;
15'b0000100111011000111 : color = 12'he73;
15'b0000100111011001000 : color = 12'he73;
15'b0000100111011001001 : color = 12'he73;
15'b0000100111011001010 : color = 12'he73;
15'b0000100111011001011 : color = 12'he73;
15'b0000100111011001100 : color = 12'he73;
15'b0000100111011001101 : color = 12'he73;
15'b0000100111011001110 : color = 12'he73;
15'b0000100111011001111 : color = 12'he73;
15'b0000100111011010000 : color = 12'he73;
15'b0000100111011010001 : color = 12'he73;
15'b0000100111011010010 : color = 12'he73;
15'b0000100111011010011 : color = 12'he73;
15'b0000100111011010100 : color = 12'he73;
15'b0000100111011010101 : color = 12'he73;
15'b0000100111011010110 : color = 12'he73;
15'b0000100111011010111 : color = 12'he73;
15'b0000100111011011000 : color = 12'he73;
15'b0000100111011011001 : color = 12'he73;
15'b0000100111011011010 : color = 12'he73;
15'b0000100111011011011 : color = 12'he73;
15'b0000100111011011100 : color = 12'he73;
15'b0000100111011011101 : color = 12'he73;
15'b0000100111011011110 : color = 12'he73;
15'b0000100111011011111 : color = 12'he73;
15'b0000100111011100000 : color = 12'he73;
15'b0000100111011100001 : color = 12'he73;
15'b0000100111011100010 : color = 12'he73;
15'b0000100111011100011 : color = 12'he73;
15'b0000100111011100100 : color = 12'he73;
15'b0000100111011100101 : color = 12'he73;
15'b0000100111011100110 : color = 12'he73;
15'b0000100111011100111 : color = 12'he73;
15'b0000100111011101000 : color = 12'he73;
15'b0000100111011101001 : color = 12'he73;
15'b0000100111011101010 : color = 12'he73;
15'b0000100111011101011 : color = 12'he73;
15'b0000100111011101100 : color = 12'he73;
15'b0000100111011101101 : color = 12'he73;
15'b0000100111011101110 : color = 12'he73;
15'b0000100111011101111 : color = 12'he73;
15'b0000100111011110000 : color = 12'he73;
15'b0000100111011110001 : color = 12'he73;
15'b0000100111011110010 : color = 12'he73;
15'b0000100111011110011 : color = 12'he73;
15'b0000100111011110100 : color = 12'he73;
15'b0000100111011110101 : color = 12'he73;
15'b0000100111011110110 : color = 12'he73;
15'b0000100111011110111 : color = 12'he73;
15'b0000100111011111000 : color = 12'he73;
15'b0000100111011111001 : color = 12'he73;
15'b0000100111011111010 : color = 12'he73;
15'b0000100111011111011 : color = 12'he73;
15'b0000100111011111100 : color = 12'he73;
15'b0000100111011111101 : color = 12'he73;
15'b0000100111011111110 : color = 12'he73;
15'b0000100111011111111 : color = 12'he73;
15'b0000100111100000000 : color = 12'he73;
15'b0000100111100000001 : color = 12'he73;
15'b0000100111100000010 : color = 12'he73;
15'b0000100111100000011 : color = 12'he73;
15'b0000100111100000100 : color = 12'he73;
15'b0000100111100000101 : color = 12'he73;
15'b0000100111100000110 : color = 12'he73;
15'b0000100111100000111 : color = 12'he73;
15'b0000100111100001000 : color = 12'he73;
15'b0000100111100001001 : color = 12'he73;
15'b0000100111100001010 : color = 12'he73;
15'b0000100111100001011 : color = 12'he73;
15'b0000100111100001100 : color = 12'he73;
15'b0000100111100001101 : color = 12'he73;
15'b0000100111100001110 : color = 12'he73;
15'b0000100111100001111 : color = 12'he73;
15'b0000100111100010000 : color = 12'he73;
15'b0000100111100010001 : color = 12'he73;
15'b0000100111100010010 : color = 12'he73;
15'b0000100111100010011 : color = 12'he73;
15'b0000100111100010100 : color = 12'he73;
15'b0000100111100010101 : color = 12'he73;
15'b0000100111100010110 : color = 12'he73;
15'b0000100111100010111 : color = 12'he73;
15'b0000100111100011000 : color = 12'he73;
15'b0000100111100011001 : color = 12'he73;
15'b0000100111100011010 : color = 12'he73;
15'b0000100111100011011 : color = 12'he73;
15'b0000100111100011100 : color = 12'he73;
15'b0000100111100011101 : color = 12'he73;
15'b0000100111100011110 : color = 12'he73;
15'b0000100111100011111 : color = 12'he73;
15'b0000100111100100000 : color = 12'he73;
15'b0000100111100100001 : color = 12'he73;
15'b0000100111100100010 : color = 12'he73;
15'b0000100111100100011 : color = 12'he73;
15'b0000100111100100100 : color = 12'he73;
15'b0000100111100100101 : color = 12'he73;
15'b0000100111100100110 : color = 12'he73;
15'b0000100111100100111 : color = 12'he73;
15'b0000100111100101000 : color = 12'he73;
15'b0000100111100101001 : color = 12'he73;
15'b0000100111100101010 : color = 12'he73;
15'b0000100111100101011 : color = 12'he73;
15'b0000100111100101100 : color = 12'he73;
15'b0000100111100101101 : color = 12'he73;
15'b0000100111100101110 : color = 12'he73;
15'b0000100111100101111 : color = 12'he73;
15'b0000100111100110000 : color = 12'he73;
15'b0000100111100110001 : color = 12'he73;
15'b0000100111100110010 : color = 12'he73;
15'b0000100111100110011 : color = 12'he73;
15'b0000100111100110100 : color = 12'he73;
15'b0000100111100110101 : color = 12'he73;
15'b0000100111100110110 : color = 12'he73;
15'b0000100111100110111 : color = 12'he73;
15'b0000100111100111000 : color = 12'he73;
15'b0000100111100111001 : color = 12'he73;
15'b0000100111100111010 : color = 12'he73;
15'b0000100111100111011 : color = 12'he73;
15'b0000100111100111100 : color = 12'he73;
15'b0000100111100111101 : color = 12'he73;
15'b0000100111100111110 : color = 12'he73;
15'b0000100111100111111 : color = 12'he73;
15'b0000100111101000000 : color = 12'he73;
15'b0000100111101000001 : color = 12'he73;
15'b0000100111101000010 : color = 12'he73;
15'b0000100111101000011 : color = 12'he73;
15'b0000100111101000100 : color = 12'he73;
15'b0000100111101000101 : color = 12'he73;
15'b0000100111101000110 : color = 12'he73;
15'b0000100111101000111 : color = 12'he73;
15'b0000100111101001000 : color = 12'he73;
15'b0000100111101001001 : color = 12'he73;
15'b0000100111101001010 : color = 12'he73;
15'b0000100111101001011 : color = 12'he73;
15'b0000100111101001100 : color = 12'he73;
15'b0000100111101001101 : color = 12'he73;
15'b0000100111101001110 : color = 12'he73;
15'b0000100111101001111 : color = 12'he73;
15'b0000100111101010000 : color = 12'he73;
15'b0000100111101010001 : color = 12'he73;
15'b0000100111101010010 : color = 12'he73;
15'b0000100111101010011 : color = 12'he73;
15'b0000100111101010100 : color = 12'he73;
15'b0000100111101010101 : color = 12'he73;
15'b0000100111101010110 : color = 12'he73;
15'b0000100111101010111 : color = 12'he73;
15'b0000100111101011000 : color = 12'he73;
15'b0000100111101011001 : color = 12'he73;
15'b0000100111101011010 : color = 12'he73;
15'b0000100111101011011 : color = 12'he73;
15'b0000100111101011100 : color = 12'he73;
15'b0000100111101011101 : color = 12'he73;
15'b0000100111101011110 : color = 12'he73;
15'b0000100111101011111 : color = 12'he73;
15'b0000100111101100000 : color = 12'he73;
15'b0000100111101100001 : color = 12'he73;
15'b0000100111101100010 : color = 12'he73;
15'b0000100111101100011 : color = 12'he73;
15'b0000100111101100100 : color = 12'he73;
15'b0000100111101100101 : color = 12'he73;
15'b0000100111101100110 : color = 12'he73;
15'b0000100111101100111 : color = 12'he73;
15'b0000100111101101000 : color = 12'he73;
15'b0000100111101101001 : color = 12'he73;
15'b0000100111101101010 : color = 12'he73;
15'b0000100111101101011 : color = 12'he73;
15'b0000100111101101100 : color = 12'he73;
15'b0000100111101101101 : color = 12'he73;
15'b0000100111101101110 : color = 12'he73;
15'b0000100111101101111 : color = 12'he73;
15'b0000100111101110000 : color = 12'he73;
15'b0000100111101110001 : color = 12'he73;
15'b0000100111101110010 : color = 12'he73;
15'b0000100111101110011 : color = 12'he73;
15'b0000100111101110100 : color = 12'he73;
15'b0000100111101110101 : color = 12'he73;
15'b0000100111101110110 : color = 12'he73;
15'b0000100111101110111 : color = 12'he73;
15'b0000100111101111000 : color = 12'he73;
15'b0000100111101111001 : color = 12'he73;
15'b0000100111101111010 : color = 12'he73;
15'b0000100111101111011 : color = 12'he73;
15'b0000100111101111100 : color = 12'he73;
15'b0000100111101111101 : color = 12'he73;
15'b0000100111101111110 : color = 12'he73;
15'b0000100111101111111 : color = 12'he73;
15'b0000100111110000000 : color = 12'he73;
15'b0000100111110000001 : color = 12'he73;
15'b0000100111110000010 : color = 12'he73;
15'b0000100111110000011 : color = 12'he73;
15'b0000100111110000100 : color = 12'he73;
15'b0000100111110000101 : color = 12'he73;
15'b0000100111110000110 : color = 12'he73;
15'b0000100111110000111 : color = 12'he73;
15'b0000100111110001000 : color = 12'he73;
15'b0000100111110001001 : color = 12'he73;
15'b0000100111110001010 : color = 12'he73;
15'b0000100111110001011 : color = 12'he73;
15'b0000100111110001100 : color = 12'he73;
15'b0000100111110001101 : color = 12'he73;
15'b0000100111110001110 : color = 12'he73;
15'b0000100111110001111 : color = 12'he73;
15'b0000100111110010000 : color = 12'he73;
15'b0000100111110010001 : color = 12'he73;
15'b0000100111110010010 : color = 12'he73;
15'b0000100111110010011 : color = 12'he73;
15'b0000100111110010100 : color = 12'he73;
15'b0000100111110010101 : color = 12'he73;
15'b0000100111110010110 : color = 12'he73;
15'b0000100111110010111 : color = 12'he73;
15'b0000100111110011000 : color = 12'he73;
15'b0000100111110011001 : color = 12'he73;
15'b0000100111110011010 : color = 12'he73;
15'b0000100111110011011 : color = 12'he73;
15'b0000100111110011100 : color = 12'he73;
15'b0000100111110011101 : color = 12'he73;
15'b0000100111110011110 : color = 12'he73;
15'b0000100111110011111 : color = 12'he73;
15'b0000100111110100000 : color = 12'he73;
15'b0000100111110100001 : color = 12'he73;
15'b0000100111110100010 : color = 12'he73;
15'b0000100111110100011 : color = 12'he73;
15'b0000100111110100100 : color = 12'he73;
15'b0000100111110100101 : color = 12'he73;
15'b0000100111110100110 : color = 12'he73;
15'b0000100111110100111 : color = 12'he73;
15'b0000100111110101000 : color = 12'he73;
15'b0000100111110101001 : color = 12'he73;
15'b0000100111110101010 : color = 12'he73;
15'b0000100111110101011 : color = 12'he73;
15'b0000100111110101100 : color = 12'he73;
15'b0000100111110101101 : color = 12'he73;
15'b0000100111110101110 : color = 12'he73;
15'b0000100111110101111 : color = 12'he73;
15'b0000100111110110000 : color = 12'he73;
15'b0000100111110110001 : color = 12'he73;
15'b0000100111110110010 : color = 12'he73;
15'b0000100111110110011 : color = 12'he73;
15'b0000100111110110100 : color = 12'he73;
15'b0000100111110110101 : color = 12'he73;
15'b0000100111110110110 : color = 12'he73;
15'b0000100111110110111 : color = 12'he73;
15'b0000100111110111000 : color = 12'he73;
15'b0000100111110111001 : color = 12'he73;
15'b0000100111110111010 : color = 12'he73;
15'b0000100111110111011 : color = 12'he73;
15'b0000100111110111100 : color = 12'he73;
15'b0000100111110111101 : color = 12'he73;
15'b0000100111110111110 : color = 12'he73;
15'b0000100111110111111 : color = 12'he73;
15'b0000100111111000000 : color = 12'he73;
15'b0000100111111000001 : color = 12'he73;
15'b0000100111111000010 : color = 12'he73;
15'b0000100111111000011 : color = 12'he73;
15'b0000100111111000100 : color = 12'he73;
15'b0000100111111000101 : color = 12'he73;
15'b0000100111111000110 : color = 12'he73;
15'b0000100111111000111 : color = 12'he73;
15'b0000100111111001000 : color = 12'he73;
15'b0000100111111001001 : color = 12'he73;
15'b0000100111111001010 : color = 12'he73;
15'b0000100111111001011 : color = 12'he73;
15'b0000100111111001100 : color = 12'he73;
15'b0000100111111001101 : color = 12'he73;
15'b0000100111111001110 : color = 12'he73;
15'b0000100111111001111 : color = 12'he73;
15'b0000100111111010000 : color = 12'he73;
15'b0000100111111010001 : color = 12'he73;
15'b0000100111111010010 : color = 12'he73;
15'b0000100111111010011 : color = 12'he73;
15'b0000100111111010100 : color = 12'he73;
15'b0000100111111010101 : color = 12'he73;
15'b0000100111111010110 : color = 12'he73;
15'b0000100111111010111 : color = 12'he73;
15'b0000100111111011000 : color = 12'he73;
15'b0000100111111011001 : color = 12'he73;
15'b0000100111111011010 : color = 12'he73;
15'b0000100111111011011 : color = 12'he73;
15'b0000100111111011100 : color = 12'he73;
15'b0000100111111011101 : color = 12'he73;
15'b0000100111111011110 : color = 12'he73;
15'b0000100111111011111 : color = 12'he73;
15'b0000100111111100000 : color = 12'he73;
15'b0000100111111100001 : color = 12'he73;
15'b0000100111111100010 : color = 12'he73;
15'b0000100111111100011 : color = 12'he73;
15'b0000100111111100100 : color = 12'he73;
15'b0000100111111100101 : color = 12'he73;
15'b0000100111111100110 : color = 12'he73;
15'b0000100111111100111 : color = 12'he73;
15'b0000100111111101000 : color = 12'he73;
15'b0000100111111101001 : color = 12'he73;
15'b0000100111111101010 : color = 12'he73;
15'b0000100111111101011 : color = 12'he73;
15'b0000100111111101100 : color = 12'he73;
15'b0000100111111101101 : color = 12'he73;
15'b0000100111111101110 : color = 12'he73;
15'b0000100111111101111 : color = 12'he73;
15'b0000100111111110000 : color = 12'he73;
15'b0000100111111110001 : color = 12'he73;
15'b0000100111111110010 : color = 12'he73;
15'b0000100111111110011 : color = 12'he73;
15'b0000100111111110100 : color = 12'he73;
15'b0000100111111110101 : color = 12'he73;
15'b0000100111111110110 : color = 12'he73;
15'b0000100111111110111 : color = 12'he73;
15'b0000100111111111000 : color = 12'he73;
15'b0000100111111111001 : color = 12'he73;
15'b0000100111111111010 : color = 12'he73;
15'b0000100111111111011 : color = 12'he73;
15'b0000100111111111100 : color = 12'he73;
15'b0000100111111111101 : color = 12'he73;
15'b0000100111111111110 : color = 12'he73;
15'b0000100111111111111 : color = 12'he73;
15'b0000101000000000000 : color = 12'he73;
15'b0000101000000000001 : color = 12'he73;
15'b0000101000000000010 : color = 12'he73;
15'b0000101000000000011 : color = 12'he73;
15'b0000101000000000100 : color = 12'he73;
15'b0000101000000000101 : color = 12'he73;
15'b0000101000000000110 : color = 12'he73;
15'b0000101000000000111 : color = 12'he73;
15'b0000101000000001000 : color = 12'he73;
15'b0000101000000001001 : color = 12'he73;
15'b0000101000000001010 : color = 12'he73;
15'b0000101000000001011 : color = 12'he73;
15'b0000101000000001100 : color = 12'he73;
15'b0000101000000001101 : color = 12'he73;
15'b0000101000000001110 : color = 12'he73;
15'b0000101000000001111 : color = 12'he73;
15'b0000101000000010000 : color = 12'he73;
15'b0000101000000010001 : color = 12'he73;
15'b0000101000000010010 : color = 12'he73;
15'b0000101000000010011 : color = 12'he73;
15'b0000101000000010100 : color = 12'he73;
15'b0000101000000010101 : color = 12'he73;
15'b0000101000000010110 : color = 12'he73;
15'b0000101000000010111 : color = 12'he73;
15'b0000101000000011000 : color = 12'he73;
15'b0000101000000011001 : color = 12'he73;
15'b0000101000000011010 : color = 12'he73;
15'b0000101000000011011 : color = 12'he73;
15'b0000101000000011100 : color = 12'he73;
15'b0000101000000011101 : color = 12'he73;
15'b0000101000000011110 : color = 12'he73;
15'b0000101000000011111 : color = 12'he73;
15'b0000101000000100000 : color = 12'he73;
15'b0000101000000100001 : color = 12'he73;
15'b0000101000000100010 : color = 12'he73;
15'b0000101000000100011 : color = 12'he73;
15'b0000101000000100100 : color = 12'he73;
15'b0000101000000100101 : color = 12'he73;
15'b0000101000000100110 : color = 12'he73;
15'b0000101000000100111 : color = 12'he73;
15'b0000101000000101000 : color = 12'he73;
15'b0000101000000101001 : color = 12'he73;
15'b0000101000000101010 : color = 12'he73;
15'b0000101000000101011 : color = 12'he73;
15'b0000101000000101100 : color = 12'he73;
15'b0000101000000101101 : color = 12'he73;
15'b0000101000000101110 : color = 12'he73;
15'b0000101000000101111 : color = 12'he73;
15'b0000101000000110000 : color = 12'he73;
15'b0000101000000110001 : color = 12'he73;
15'b0000101000000110010 : color = 12'he73;
15'b0000101000000110011 : color = 12'he73;
15'b0000101000000110100 : color = 12'he73;
15'b0000101000000110101 : color = 12'he73;
15'b0000101000000110110 : color = 12'he73;
15'b0000101000000110111 : color = 12'he73;
15'b0000101000000111000 : color = 12'he73;
15'b0000101000000111001 : color = 12'he73;
15'b0000101000000111010 : color = 12'he73;
15'b0000101000000111011 : color = 12'he73;
15'b0000101000000111100 : color = 12'he73;
15'b0000101000000111101 : color = 12'he73;
15'b0000101000000111110 : color = 12'he73;
15'b0000101000000111111 : color = 12'he73;
15'b0000101000001000000 : color = 12'he73;
15'b0000101000001000001 : color = 12'he73;
15'b0000101000001000010 : color = 12'he73;
15'b0000101000001000011 : color = 12'he73;
15'b0000101000001000100 : color = 12'he73;
15'b0000101000001000101 : color = 12'he73;
15'b0000101000001000110 : color = 12'he73;
15'b0000101000001000111 : color = 12'he73;
15'b0000101000001001000 : color = 12'he73;
15'b0000101000001001001 : color = 12'he73;
15'b0000101000001001010 : color = 12'he73;
15'b0000101000001001011 : color = 12'he73;
15'b0000101000001001100 : color = 12'he73;
15'b0000101000001001101 : color = 12'he73;
15'b0000101000001001110 : color = 12'he73;
15'b0000101000001001111 : color = 12'he73;
15'b0000101000001010000 : color = 12'he73;
15'b0000101000001010001 : color = 12'he73;
15'b0000101000001010010 : color = 12'he73;
15'b0000101000001010011 : color = 12'he73;
15'b0000101000001010100 : color = 12'he73;
15'b0000101000001010101 : color = 12'he73;
15'b0000101000001010110 : color = 12'he73;
15'b0000101000001010111 : color = 12'he73;
15'b0000101000001011000 : color = 12'he73;
15'b0000101000001011001 : color = 12'he73;
15'b0000101000001011010 : color = 12'he73;
15'b0000101000001011011 : color = 12'he73;
15'b0000101000001011100 : color = 12'he73;
15'b0000101000001011101 : color = 12'he73;
15'b0000101000001011110 : color = 12'he73;
15'b0000101000001011111 : color = 12'he73;
15'b0000101000001100000 : color = 12'he73;
15'b0000101000001100001 : color = 12'he73;
15'b0000101000001100010 : color = 12'he73;
15'b0000101000001100011 : color = 12'he73;
15'b0000101000001100100 : color = 12'he73;
15'b0000101000001100101 : color = 12'he73;
15'b0000101000001100110 : color = 12'he73;
15'b0000101000001100111 : color = 12'he73;
15'b0000101000001101000 : color = 12'he73;
15'b0000101000001101001 : color = 12'he73;
15'b0000101000001101010 : color = 12'he73;
15'b0000101000001101011 : color = 12'he73;
15'b0000101000001101100 : color = 12'he73;
15'b0000101000001101101 : color = 12'he73;
15'b0000101000001101110 : color = 12'he73;
15'b0000101000001101111 : color = 12'he73;
15'b0000101000001110000 : color = 12'he73;
15'b0000101000001110001 : color = 12'he73;
15'b0000101000001110010 : color = 12'he73;
15'b0000101000001110011 : color = 12'he73;
15'b0000101000001110100 : color = 12'he73;
15'b0000101000001110101 : color = 12'he73;
15'b0000101000001110110 : color = 12'he73;
15'b0000101000001110111 : color = 12'he73;
15'b0000101000001111000 : color = 12'he73;
15'b0000101000001111001 : color = 12'he73;
15'b0000101000001111010 : color = 12'he73;
15'b0000101000001111011 : color = 12'he73;
15'b0000101000001111100 : color = 12'he73;
15'b0000101000001111101 : color = 12'he73;
15'b0000101000001111110 : color = 12'he73;
15'b0000101000001111111 : color = 12'he73;
15'b0000101000010000000 : color = 12'he73;
15'b0000101000010000001 : color = 12'he73;
15'b0000101000010000010 : color = 12'he73;
15'b0000101000010000011 : color = 12'he73;
15'b0000101000010000100 : color = 12'he73;
15'b0000101000010000101 : color = 12'he73;
15'b0000101000010000110 : color = 12'he73;
15'b0000101000010000111 : color = 12'he73;
15'b0000101000010001000 : color = 12'he73;
15'b0000101000010001001 : color = 12'he73;
15'b0000101000010001010 : color = 12'he73;
15'b0000101000010001011 : color = 12'he73;
15'b0000101000010001100 : color = 12'he73;
15'b0000101000010001101 : color = 12'he73;
15'b0000100111011001100 : color = 12'he73;
15'b0000100111011001101 : color = 12'he73;
15'b0000100111011001110 : color = 12'he73;
15'b0000100111011001111 : color = 12'he73;
15'b0000100111011010000 : color = 12'he73;
15'b0000100111011010001 : color = 12'he73;
15'b0000100111011010010 : color = 12'he73;
15'b0000100111011010011 : color = 12'he73;
15'b0000100111011010100 : color = 12'he73;
15'b0000100111011010101 : color = 12'he73;
15'b0000100111011010110 : color = 12'he73;
15'b0000100111011010111 : color = 12'he73;
15'b0000100111011011000 : color = 12'he73;
15'b0000100111011011001 : color = 12'he73;
15'b0000100111011011010 : color = 12'he73;
15'b0000100111011011011 : color = 12'he73;
15'b0000100111011011100 : color = 12'he73;
15'b0000100111011011101 : color = 12'he73;
15'b0000100111011011110 : color = 12'he73;
15'b0000100111011011111 : color = 12'he73;
15'b0000100111011100000 : color = 12'he73;
15'b0000100111011100001 : color = 12'he73;
15'b0000100111011100010 : color = 12'he73;
15'b0000100111011100011 : color = 12'he73;
15'b0000100111011100100 : color = 12'he73;
15'b0000100111011100101 : color = 12'he73;
15'b0000100111011100110 : color = 12'he73;
15'b0000100111011100111 : color = 12'he73;
15'b0000100111011101000 : color = 12'he73;
15'b0000100111011101001 : color = 12'he73;
15'b0000100111011101010 : color = 12'he73;
15'b0000100111011101011 : color = 12'he73;
15'b0000100111011101100 : color = 12'he73;
15'b0000100111011101101 : color = 12'he73;
15'b0000100111011101110 : color = 12'he73;
15'b0000100111011101111 : color = 12'he73;
15'b0000100111011110000 : color = 12'he73;
15'b0000100111011110001 : color = 12'he73;
15'b0000100111011110010 : color = 12'he73;
15'b0000100111011110011 : color = 12'he73;
15'b0000100111011110100 : color = 12'he73;
15'b0000100111011110101 : color = 12'he73;
15'b0000100111011110110 : color = 12'he73;
15'b0000100111011110111 : color = 12'he73;
15'b0000100111011111000 : color = 12'he73;
15'b0000100111011111001 : color = 12'he73;
15'b0000100111011111010 : color = 12'he73;
15'b0000100111011111011 : color = 12'he73;
15'b0000100111011111100 : color = 12'he73;
15'b0000100111011111101 : color = 12'he73;
15'b0000100111011111110 : color = 12'he73;
15'b0000100111011111111 : color = 12'he73;
15'b0000100111100000000 : color = 12'he73;
15'b0000100111100000001 : color = 12'he73;
15'b0000100111100000010 : color = 12'he73;
15'b0000100111100000011 : color = 12'he73;
15'b0000100111100000100 : color = 12'he73;
15'b0000100111100000101 : color = 12'he73;
15'b0000100111100000110 : color = 12'he73;
15'b0000100111100000111 : color = 12'he73;
15'b0000100111100001000 : color = 12'he73;
15'b0000100111100001001 : color = 12'he73;
15'b0000100111100001010 : color = 12'he73;
15'b0000100111100001011 : color = 12'he73;
15'b0000100111100001100 : color = 12'he73;
15'b0000100111100001101 : color = 12'he73;
15'b0000100111100001110 : color = 12'he73;
15'b0000100111100001111 : color = 12'he73;
15'b0000100111100010000 : color = 12'he73;
15'b0000100111100010001 : color = 12'he73;
15'b0000100111100010010 : color = 12'he73;
15'b0000100111100010011 : color = 12'he73;
15'b0000100111100010100 : color = 12'he73;
15'b0000100111100010101 : color = 12'he73;
15'b0000100111100010110 : color = 12'he73;
15'b0000100111100010111 : color = 12'he73;
15'b0000100111100011000 : color = 12'he73;
15'b0000100111100011001 : color = 12'he73;
15'b0000100111100011010 : color = 12'he73;
15'b0000100111100011011 : color = 12'he73;
15'b0000100111100011100 : color = 12'he73;
15'b0000100111100011101 : color = 12'he73;
15'b0000100111100011110 : color = 12'he73;
15'b0000100111100011111 : color = 12'he73;
15'b0000100111100100000 : color = 12'he73;
15'b0000100111100100001 : color = 12'he73;
15'b0000100111100100010 : color = 12'he73;
15'b0000100111100100011 : color = 12'he73;
15'b0000100111100100100 : color = 12'he73;
15'b0000100111100100101 : color = 12'he73;
15'b0000100111100100110 : color = 12'he73;
15'b0000100111100100111 : color = 12'he73;
15'b0000100111100101000 : color = 12'he73;
15'b0000100111100101001 : color = 12'he73;
15'b0000100111100101010 : color = 12'he73;
15'b0000100111100101011 : color = 12'he73;
15'b0000100111100101100 : color = 12'he73;
15'b0000100111100101101 : color = 12'he73;
15'b0000100111100101110 : color = 12'he73;
15'b0000100111100101111 : color = 12'he73;
15'b0000100111100110000 : color = 12'he73;
15'b0000100111100110001 : color = 12'he73;
15'b0000100111100110010 : color = 12'he73;
15'b0000100111100110011 : color = 12'he73;
15'b0000100111100110100 : color = 12'he73;
15'b0000100111100110101 : color = 12'he73;
15'b0000100111100110110 : color = 12'he73;
15'b0000100111100110111 : color = 12'he73;
15'b0000100111100111000 : color = 12'he73;
15'b0000100111100111001 : color = 12'he73;
15'b0000100111100111010 : color = 12'he73;
15'b0000100111100111011 : color = 12'he73;
15'b0000100111100111100 : color = 12'he73;
15'b0000100111100111101 : color = 12'he73;
15'b0000100111100111110 : color = 12'he73;
15'b0000100111100111111 : color = 12'he73;
15'b0000100111101000000 : color = 12'he73;
15'b0000100111101000001 : color = 12'he73;
15'b0000100111101000010 : color = 12'he73;
15'b0000100111101000011 : color = 12'he73;
15'b0000100111101000100 : color = 12'he73;
15'b0000100111101000101 : color = 12'he73;
15'b0000100111101000110 : color = 12'he73;
15'b0000100111101000111 : color = 12'he73;
15'b0000100111101001000 : color = 12'he73;
15'b0000100111101001001 : color = 12'he73;
15'b0000100111101001010 : color = 12'he73;
15'b0000100111101001011 : color = 12'he73;
15'b0000100111101001100 : color = 12'he73;
15'b0000100111101001101 : color = 12'he73;
15'b0000100111101001110 : color = 12'he73;
15'b0000100111101001111 : color = 12'he73;
15'b0000100111101010000 : color = 12'he73;
15'b0000100111101010001 : color = 12'he73;
15'b0000100111101010010 : color = 12'he73;
15'b0000100111101010011 : color = 12'he73;
15'b0000100111101010100 : color = 12'he73;
15'b0000100111101010101 : color = 12'he73;
15'b0000100111101010110 : color = 12'he73;
15'b0000100111101010111 : color = 12'he73;
15'b0000100111101011000 : color = 12'he73;
15'b0000100111101011001 : color = 12'he73;
15'b0000100111101011010 : color = 12'he73;
15'b0000100111101011011 : color = 12'he73;
15'b0000100111101011100 : color = 12'he73;
15'b0000100111101011101 : color = 12'he73;
15'b0000100111101011110 : color = 12'he73;
15'b0000100111101011111 : color = 12'he73;
15'b0000100111101100000 : color = 12'he73;
15'b0000100111101100001 : color = 12'he73;
15'b0000100111101100010 : color = 12'he73;
15'b0000100111101100011 : color = 12'he73;
15'b0000100111101100100 : color = 12'he73;
15'b0000100111101100101 : color = 12'he73;
15'b0000100111101100110 : color = 12'he73;
15'b0000100111101100111 : color = 12'he73;
15'b0000100111101101000 : color = 12'he73;
15'b0000100111101101001 : color = 12'he73;
15'b0000100111101101010 : color = 12'he73;
15'b0000100111101101011 : color = 12'he73;
15'b0000100111101101100 : color = 12'he73;
15'b0000100111101101101 : color = 12'he73;
15'b0000100111101101110 : color = 12'he73;
15'b0000100111101101111 : color = 12'he73;
15'b0000100111101110000 : color = 12'he73;
15'b0000100111101110001 : color = 12'he73;
15'b0000100111101110010 : color = 12'he73;
15'b0000100111101110011 : color = 12'he73;
15'b0000100111101110100 : color = 12'he73;
15'b0000100111101110101 : color = 12'he73;
15'b0000100111101110110 : color = 12'he73;
15'b0000100111101110111 : color = 12'he73;
15'b0000100111101111000 : color = 12'he73;
15'b0000100111101111001 : color = 12'he73;
15'b0000100111101111010 : color = 12'he73;
15'b0000100111101111011 : color = 12'he73;
15'b0000100111101111100 : color = 12'he73;
15'b0000100111101111101 : color = 12'he73;
15'b0000100111101111110 : color = 12'he73;
15'b0000100111101111111 : color = 12'he73;
15'b0000100111110000000 : color = 12'he73;
15'b0000100111110000001 : color = 12'he73;
15'b0000100111110000010 : color = 12'he73;
15'b0000100111110000011 : color = 12'he73;
15'b0000100111110000100 : color = 12'he73;
15'b0000100111110000101 : color = 12'he73;
15'b0000100111110000110 : color = 12'he73;
15'b0000100111110000111 : color = 12'he73;
15'b0000100111110001000 : color = 12'he73;
15'b0000100111110001001 : color = 12'he73;
15'b0000100111110001010 : color = 12'he73;
15'b0000100111110001011 : color = 12'he73;
15'b0000100111110001100 : color = 12'he73;
15'b0000100111110001101 : color = 12'he73;
15'b0000100111110001110 : color = 12'he73;
15'b0000100111110001111 : color = 12'he73;
15'b0000100111110010000 : color = 12'he73;
15'b0000100111110010001 : color = 12'he73;
15'b0000100111110010010 : color = 12'he73;
15'b0000100111110010011 : color = 12'he73;
15'b0000100111110010100 : color = 12'he73;
15'b0000100111110010101 : color = 12'he73;
15'b0000100111110010110 : color = 12'he73;
15'b0000100111110010111 : color = 12'he73;
15'b0000100111110011000 : color = 12'he73;
15'b0000100111110011001 : color = 12'he73;
15'b0000100111110011010 : color = 12'he73;
15'b0000100111110011011 : color = 12'he73;
15'b0000100111110011100 : color = 12'he73;
15'b0000100111110011101 : color = 12'he73;
15'b0000100111110011110 : color = 12'he73;
15'b0000100111110011111 : color = 12'he73;
15'b0000100111110100000 : color = 12'he73;
15'b0000100111110100001 : color = 12'he73;
15'b0000100111110100010 : color = 12'he73;
15'b0000100111110100011 : color = 12'he73;
15'b0000100111110100100 : color = 12'he73;
15'b0000100111110100101 : color = 12'he73;
15'b0000100111110100110 : color = 12'he73;
15'b0000100111110100111 : color = 12'he73;
15'b0000100111110101000 : color = 12'he73;
15'b0000100111110101001 : color = 12'he73;
15'b0000100111110101010 : color = 12'he73;
15'b0000100111110101011 : color = 12'he73;
15'b0000100111110101100 : color = 12'he73;
15'b0000100111110101101 : color = 12'he73;
15'b0000100111110101110 : color = 12'he73;
15'b0000100111110101111 : color = 12'he73;
15'b0000100111110110000 : color = 12'he73;
15'b0000100111110110001 : color = 12'he73;
15'b0000100111110110010 : color = 12'he73;
15'b0000100111110110011 : color = 12'he73;
15'b0000100111110110100 : color = 12'he73;
15'b0000100111110110101 : color = 12'he73;
15'b0000100111110110110 : color = 12'he73;
15'b0000100111110110111 : color = 12'he73;
15'b0000100111110111000 : color = 12'he73;
15'b0000100111110111001 : color = 12'he73;
15'b0000100111110111010 : color = 12'he73;
15'b0000100111110111011 : color = 12'he73;
15'b0000100111110111100 : color = 12'he73;
15'b0000100111110111101 : color = 12'he73;
15'b0000100111110111110 : color = 12'he73;
15'b0000100111110111111 : color = 12'he73;
15'b0000100111111000000 : color = 12'he73;
15'b0000100111111000001 : color = 12'he73;
15'b0000100111111000010 : color = 12'he73;
15'b0000100111111000011 : color = 12'he73;
15'b0000100111111000100 : color = 12'he73;
15'b0000100111111000101 : color = 12'he73;
15'b0000100111111000110 : color = 12'he73;
15'b0000100111111000111 : color = 12'he73;
15'b0000100111111001000 : color = 12'he73;
15'b0000100111111001001 : color = 12'he73;
15'b0000100111111001010 : color = 12'he73;
15'b0000100111111001011 : color = 12'he73;
15'b0000100111111001100 : color = 12'he73;
15'b0000100111111001101 : color = 12'he73;
15'b0000100111111001110 : color = 12'he73;
15'b0000100111111001111 : color = 12'he73;
15'b0000100111111010000 : color = 12'he73;
15'b0000100111111010001 : color = 12'he73;
15'b0000100111111010010 : color = 12'he73;
15'b0000100111111010011 : color = 12'he73;
15'b0000100111111010100 : color = 12'he73;
15'b0000100111111010101 : color = 12'he73;
15'b0000100111111010110 : color = 12'he73;
15'b0000100111111010111 : color = 12'he73;
15'b0000100111111011000 : color = 12'he73;
15'b0000100111111011001 : color = 12'he73;
15'b0000100111111011010 : color = 12'he73;
15'b0000100111111011011 : color = 12'he73;
15'b0000100111111011100 : color = 12'he73;
15'b0000100111111011101 : color = 12'he73;
15'b0000100111111011110 : color = 12'he73;
15'b0000100111111011111 : color = 12'he73;
15'b0000100111111100000 : color = 12'he73;
15'b0000100111111100001 : color = 12'he73;
15'b0000100111111100010 : color = 12'he73;
15'b0000100111111100011 : color = 12'he73;
15'b0000100111111100100 : color = 12'he73;
15'b0000100111111100101 : color = 12'he73;
15'b0000100111111100110 : color = 12'he73;
15'b0000100111111100111 : color = 12'he73;
15'b0000100111111101000 : color = 12'he73;
15'b0000100111111101001 : color = 12'he73;
15'b0000100111111101010 : color = 12'he73;
15'b0000100111111101011 : color = 12'he73;
15'b0000100111111101100 : color = 12'he73;
15'b0000100111111101101 : color = 12'he73;
15'b0000100111111101110 : color = 12'he73;
15'b0000100111111101111 : color = 12'he73;
15'b0000100111111110000 : color = 12'he73;
15'b0000100111111110001 : color = 12'he73;
15'b0000100111111110010 : color = 12'he73;
15'b0000100111111110011 : color = 12'he73;
15'b0000100111111110100 : color = 12'he73;
15'b0000100111111110101 : color = 12'he73;
15'b0000100111111110110 : color = 12'he73;
15'b0000100111111110111 : color = 12'he73;
15'b0000100111111111000 : color = 12'he73;
15'b0000100111111111001 : color = 12'he73;
15'b0000100111111111010 : color = 12'he73;
15'b0000100111111111011 : color = 12'he73;
15'b0000100111111111100 : color = 12'he73;
15'b0000100111111111101 : color = 12'he73;
15'b0000100111111111110 : color = 12'he73;
15'b0000100111111111111 : color = 12'he73;
15'b0000101000000000000 : color = 12'he73;
15'b0000101000000000001 : color = 12'he73;
15'b0000101000000000010 : color = 12'he73;
15'b0000101000000000011 : color = 12'he73;
15'b0000101000000000100 : color = 12'he73;
15'b0000101000000000101 : color = 12'he73;
15'b0000101000000000110 : color = 12'he73;
15'b0000101000000000111 : color = 12'he73;
15'b0000101000000001000 : color = 12'he73;
15'b0000101000000001001 : color = 12'he73;
15'b0000101000000001010 : color = 12'he73;
15'b0000101000000001011 : color = 12'he73;
15'b0000101000000001100 : color = 12'he73;
15'b0000101000000001101 : color = 12'he73;
15'b0000101000000001110 : color = 12'he73;
15'b0000101000000001111 : color = 12'he73;
15'b0000101000000010000 : color = 12'he73;
15'b0000101000000010001 : color = 12'he73;
15'b0000101000000010010 : color = 12'he73;
15'b0000101000000010011 : color = 12'he73;
15'b0000101000000010100 : color = 12'he73;
15'b0000101000000010101 : color = 12'he73;
15'b0000101000000010110 : color = 12'he73;
15'b0000101000000010111 : color = 12'he73;
15'b0000101000000011000 : color = 12'he73;
15'b0000101000000011001 : color = 12'he73;
15'b0000101000000011010 : color = 12'he73;
15'b0000101000000011011 : color = 12'he73;
15'b0000101000000011100 : color = 12'he73;
15'b0000101000000011101 : color = 12'he73;
15'b0000101000000011110 : color = 12'he73;
15'b0000101000000011111 : color = 12'he73;
15'b0000101000000100000 : color = 12'he73;
15'b0000101000000100001 : color = 12'he73;
15'b0000101000000100010 : color = 12'he73;
15'b0000101000000100011 : color = 12'he73;
15'b0000101000000100100 : color = 12'he73;
15'b0000101000000100101 : color = 12'he73;
15'b0000101000000100110 : color = 12'he73;
15'b0000101000000100111 : color = 12'he73;
15'b0000101000000101000 : color = 12'he73;
15'b0000101000000101001 : color = 12'he73;
15'b0000101000000101010 : color = 12'he73;
15'b0000101000000101011 : color = 12'he73;
15'b0000101000000101100 : color = 12'he73;
15'b0000101000000101101 : color = 12'he73;
15'b0000101000000101110 : color = 12'he73;
15'b0000101000000101111 : color = 12'he73;
15'b0000101000000110000 : color = 12'he73;
15'b0000101000000110001 : color = 12'he73;
15'b0000101000000110010 : color = 12'he73;
15'b0000101000000110011 : color = 12'he73;
15'b0000101000000110100 : color = 12'he73;
15'b0000101000000110101 : color = 12'he73;
15'b0000101000000110110 : color = 12'he73;
15'b0000101000000110111 : color = 12'he73;
15'b0000101000000111000 : color = 12'he73;
15'b0000101000000111001 : color = 12'he73;
15'b0000101000000111010 : color = 12'he73;
15'b0000101000000111011 : color = 12'he73;
15'b0000101000000111100 : color = 12'he73;
15'b0000101000000111101 : color = 12'he73;
15'b0000101000000111110 : color = 12'he73;
15'b0000101000000111111 : color = 12'he73;
15'b0000101000001000000 : color = 12'he73;
15'b0000101000001000001 : color = 12'he73;
15'b0000101000001000010 : color = 12'he73;
15'b0000101000001000011 : color = 12'he73;
15'b0000101000001000100 : color = 12'he73;
15'b0000101000001000101 : color = 12'he73;
15'b0000101000001000110 : color = 12'he73;
15'b0000101000001000111 : color = 12'he73;
15'b0000101000001001000 : color = 12'he73;
15'b0000101000001001001 : color = 12'he73;
15'b0000101000001001010 : color = 12'he73;
15'b0000101000001001011 : color = 12'he73;
15'b0000101000001001100 : color = 12'he73;
15'b0000101000001001101 : color = 12'he73;
15'b0000101000001001110 : color = 12'he73;
15'b0000101000001001111 : color = 12'he73;
15'b0000101000001010000 : color = 12'he73;
15'b0000101000001010001 : color = 12'he73;
15'b0000101000001010010 : color = 12'he73;
15'b0000101000001010011 : color = 12'he73;
15'b0000101000001010100 : color = 12'he73;
15'b0000101000001010101 : color = 12'he73;
15'b0000101000001010110 : color = 12'he73;
15'b0000101000001010111 : color = 12'he73;
15'b0000101000001011000 : color = 12'he73;
15'b0000101000001011001 : color = 12'he73;
15'b0000101000001011010 : color = 12'he73;
15'b0000101000001011011 : color = 12'he73;
15'b0000101000001011100 : color = 12'he73;
15'b0000101000001011101 : color = 12'he73;
15'b0000101000001011110 : color = 12'he73;
15'b0000101000001011111 : color = 12'he73;
15'b0000101000001100000 : color = 12'he73;
15'b0000101000001100001 : color = 12'he73;
15'b0000101000001100010 : color = 12'he73;
15'b0000101000001100011 : color = 12'he73;
15'b0000101000001100100 : color = 12'he73;
15'b0000101000001100101 : color = 12'he73;
15'b0000101000001100110 : color = 12'he73;
15'b0000101000001100111 : color = 12'he73;
15'b0000101000001101000 : color = 12'he73;
15'b0000101000001101001 : color = 12'he73;
15'b0000101000001101010 : color = 12'he73;
15'b0000101000001101011 : color = 12'he73;
15'b0000101000001101100 : color = 12'he73;
15'b0000101000001101101 : color = 12'he73;
15'b0000101000001101110 : color = 12'he73;
15'b0000101000001101111 : color = 12'he73;
15'b0000101000001110000 : color = 12'he73;
15'b0000101000001110001 : color = 12'he73;
15'b0000101000001110010 : color = 12'he73;
15'b0000101000001110011 : color = 12'he73;
15'b0000101000001110100 : color = 12'he73;
15'b0000101000001110101 : color = 12'he73;
15'b0000101000001110110 : color = 12'he73;
15'b0000101000001110111 : color = 12'he73;
15'b0000101000001111000 : color = 12'he73;
15'b0000101000001111001 : color = 12'he73;
15'b0000101000001111010 : color = 12'he73;
15'b0000101000001111011 : color = 12'he73;
15'b0000101000001111100 : color = 12'he73;
15'b0000101000001111101 : color = 12'he73;
15'b0000101000001111110 : color = 12'he73;
15'b0000101000001111111 : color = 12'he73;
15'b0000101000010000000 : color = 12'he73;
15'b0000101000010000001 : color = 12'he73;
15'b0000101000010000010 : color = 12'he73;
15'b0000101000010000011 : color = 12'he73;
15'b0000101000010000100 : color = 12'he73;
15'b0000101000010000101 : color = 12'he73;
15'b0000101000010000110 : color = 12'he73;
15'b0000101000010000111 : color = 12'he73;
15'b0000101000010001000 : color = 12'he73;
15'b0000101000010001001 : color = 12'he73;
15'b0000101000010001010 : color = 12'he73;
15'b0000101000010001011 : color = 12'he73;
15'b0000101000010001100 : color = 12'he73;
15'b0000101000010001101 : color = 12'he73;
15'b0000101000010001110 : color = 12'he73;
15'b0000101000010001111 : color = 12'he73;
15'b0000101000010010000 : color = 12'he73;
15'b0000101000010010001 : color = 12'he73;
15'b0000101000010010010 : color = 12'he73;
15'b0000101000010010011 : color = 12'he73;
15'b0000101000010010100 : color = 12'he73;
15'b0000101000010010101 : color = 12'he73;
15'b0000101000010010110 : color = 12'he73;
15'b0000101000010010111 : color = 12'he73;
15'b0000101000010011000 : color = 12'he73;
15'b0000101000010011001 : color = 12'he73;
15'b0000101000010011010 : color = 12'he73;
15'b0000101000010011011 : color = 12'he73;
15'b0000101000010011100 : color = 12'he73;
15'b0000101000010011101 : color = 12'he73;
15'b0000101000010011110 : color = 12'he73;
15'b0000101000010011111 : color = 12'he73;
15'b0000101000010100000 : color = 12'he73;
15'b0000101000010100001 : color = 12'he73;
15'b0000101000010100010 : color = 12'he73;
15'b0000101000010100011 : color = 12'he73;
15'b0000101000010100100 : color = 12'he73;
15'b0000101000010100101 : color = 12'he73;
15'b0000101000010100110 : color = 12'he73;
15'b0000101000010100111 : color = 12'he73;
15'b0000101000010101000 : color = 12'he73;
15'b0000101000010101001 : color = 12'he73;
15'b0000101000010101010 : color = 12'he73;
15'b0000101000010101011 : color = 12'he73;
15'b0000101000010101100 : color = 12'he73;
15'b0000101000010101101 : color = 12'he73;
15'b0000101000010101110 : color = 12'he73;
15'b0000101000010101111 : color = 12'he73;
15'b0000101000010110000 : color = 12'he73;
15'b0000101000010110001 : color = 12'he73;
15'b0000101000010110010 : color = 12'he73;
15'b0000101000010110011 : color = 12'he73;
15'b0000101000010110100 : color = 12'he73;
15'b0000101000010110101 : color = 12'he73;
15'b0000101000010110110 : color = 12'he73;
15'b0000100111011110101 : color = 12'he73;
15'b0000100111011110110 : color = 12'he73;
15'b0000100111011110111 : color = 12'he73;
15'b0000100111011111000 : color = 12'he73;
15'b0000100111011111001 : color = 12'he73;
15'b0000100111011111010 : color = 12'he73;
15'b0000100111011111011 : color = 12'he73;
15'b0000100111011111100 : color = 12'he73;
15'b0000100111011111101 : color = 12'he73;
15'b0000100111011111110 : color = 12'he73;
15'b0000100111011111111 : color = 12'he73;
15'b0000100111100000000 : color = 12'he73;
15'b0000100111100000001 : color = 12'he73;
15'b0000100111100000010 : color = 12'he73;
15'b0000100111100000011 : color = 12'he73;
15'b0000100111100000100 : color = 12'he73;
15'b0000100111100000101 : color = 12'he73;
15'b0000100111100000110 : color = 12'he73;
15'b0000100111100000111 : color = 12'he73;
15'b0000100111100001000 : color = 12'he73;
15'b0000100111100001001 : color = 12'he73;
15'b0000100111100001010 : color = 12'he73;
15'b0000100111100001011 : color = 12'he73;
15'b0000100111100001100 : color = 12'he73;
15'b0000100111100001101 : color = 12'he73;
15'b0000100111100001110 : color = 12'he73;
15'b0000100111100001111 : color = 12'he73;
15'b0000100111100010000 : color = 12'he73;
15'b0000100111100010001 : color = 12'he73;
15'b0000100111100010010 : color = 12'he73;
15'b0000100111100010011 : color = 12'he73;
15'b0000100111100010100 : color = 12'he73;
15'b0000100111100010101 : color = 12'he73;
15'b0000100111100010110 : color = 12'he73;
15'b0000100111100010111 : color = 12'he73;
15'b0000100111100011000 : color = 12'he73;
15'b0000100111100011001 : color = 12'he73;
15'b0000100111100011010 : color = 12'he73;
15'b0000100111100011011 : color = 12'he73;
15'b0000100111100011100 : color = 12'he73;
15'b0000100111100011101 : color = 12'he73;
15'b0000100111100011110 : color = 12'he73;
15'b0000100111100011111 : color = 12'he73;
15'b0000100111100100000 : color = 12'he73;
15'b0000100111100100001 : color = 12'he73;
15'b0000100111100100010 : color = 12'he73;
15'b0000100111100100011 : color = 12'he73;
15'b0000100111100100100 : color = 12'he73;
15'b0000100111100100101 : color = 12'he73;
15'b0000100111100100110 : color = 12'he73;
15'b0000100111100100111 : color = 12'he73;
15'b0000100111100101000 : color = 12'he73;
15'b0000100111100101001 : color = 12'he73;
15'b0000100111100101010 : color = 12'he73;
15'b0000100111100101011 : color = 12'he73;
15'b0000100111100101100 : color = 12'he73;
15'b0000100111100101101 : color = 12'he73;
15'b0000100111100101110 : color = 12'he73;
15'b0000100111100101111 : color = 12'he73;
15'b0000100111100110000 : color = 12'he73;
15'b0000100111100110001 : color = 12'he73;
15'b0000100111100110010 : color = 12'he73;
15'b0000100111100110011 : color = 12'he73;
15'b0000100111100110100 : color = 12'he73;
15'b0000100111100110101 : color = 12'he73;
15'b0000100111100110110 : color = 12'he73;
15'b0000100111100110111 : color = 12'he73;
15'b0000100111100111000 : color = 12'he73;
15'b0000100111100111001 : color = 12'he73;
15'b0000100111100111010 : color = 12'he73;
15'b0000100111100111011 : color = 12'he73;
15'b0000100111100111100 : color = 12'he73;
15'b0000100111100111101 : color = 12'he73;
15'b0000100111100111110 : color = 12'he73;
15'b0000100111100111111 : color = 12'he73;
15'b0000100111101000000 : color = 12'he73;
15'b0000100111101000001 : color = 12'he73;
15'b0000100111101000010 : color = 12'he73;
15'b0000100111101000011 : color = 12'he73;
15'b0000100111101000100 : color = 12'he73;
15'b0000100111101000101 : color = 12'he73;
15'b0000100111101000110 : color = 12'he73;
15'b0000100111101000111 : color = 12'he73;
15'b0000100111101001000 : color = 12'he73;
15'b0000100111101001001 : color = 12'he73;
15'b0000100111101001010 : color = 12'he73;
15'b0000100111101001011 : color = 12'he73;
15'b0000100111101001100 : color = 12'he73;
15'b0000100111101001101 : color = 12'he73;
15'b0000100111101001110 : color = 12'he73;
15'b0000100111101001111 : color = 12'he73;
15'b0000100111101010000 : color = 12'he73;
15'b0000100111101010001 : color = 12'he73;
15'b0000100111101010010 : color = 12'he73;
15'b0000100111101010011 : color = 12'he73;
15'b0000100111101010100 : color = 12'he73;
15'b0000100111101010101 : color = 12'he73;
15'b0000100111101010110 : color = 12'he73;
15'b0000100111101010111 : color = 12'he73;
15'b0000100111101011000 : color = 12'he73;
15'b0000100111101011001 : color = 12'he73;
15'b0000100111101011010 : color = 12'he73;
15'b0000100111101011011 : color = 12'he73;
15'b0000100111101011100 : color = 12'he73;
15'b0000100111101011101 : color = 12'he73;
15'b0000100111101011110 : color = 12'he73;
15'b0000100111101011111 : color = 12'he73;
15'b0000100111101100000 : color = 12'he73;
15'b0000100111101100001 : color = 12'he73;
15'b0000100111101100010 : color = 12'he73;
15'b0000100111101100011 : color = 12'he73;
15'b0000100111101100100 : color = 12'he73;
15'b0000100111101100101 : color = 12'he73;
15'b0000100111101100110 : color = 12'he73;
15'b0000100111101100111 : color = 12'he73;
15'b0000100111101101000 : color = 12'he73;
15'b0000100111101101001 : color = 12'he73;
15'b0000100111101101010 : color = 12'he73;
15'b0000100111101101011 : color = 12'he73;
15'b0000100111101101100 : color = 12'he73;
15'b0000100111101101101 : color = 12'he73;
15'b0000100111101101110 : color = 12'he73;
15'b0000100111101101111 : color = 12'he73;
15'b0000100111101110000 : color = 12'he73;
15'b0000100111101110001 : color = 12'he73;
15'b0000100111101110010 : color = 12'he73;
15'b0000100111101110011 : color = 12'he73;
15'b0000100111101110100 : color = 12'he73;
15'b0000100111101110101 : color = 12'he73;
15'b0000100111101110110 : color = 12'he73;
15'b0000100111101110111 : color = 12'he73;
15'b0000100111101111000 : color = 12'he73;
15'b0000100111101111001 : color = 12'he73;
15'b0000100111101111010 : color = 12'he73;
15'b0000100111101111011 : color = 12'he73;
15'b0000100111101111100 : color = 12'he73;
15'b0000100111101111101 : color = 12'he73;
15'b0000100111101111110 : color = 12'he73;
15'b0000100111101111111 : color = 12'he73;
15'b0000100111110000000 : color = 12'he73;
15'b0000100111110000001 : color = 12'he73;
15'b0000100111110000010 : color = 12'he73;
15'b0000100111110000011 : color = 12'he73;
15'b0000100111110000100 : color = 12'he73;
15'b0000100111110000101 : color = 12'he73;
15'b0000100111110000110 : color = 12'he73;
15'b0000100111110000111 : color = 12'he73;
15'b0000100111110001000 : color = 12'he73;
15'b0000100111110001001 : color = 12'he73;
15'b0000100111110001010 : color = 12'he73;
15'b0000100111110001011 : color = 12'he73;
15'b0000100111110001100 : color = 12'he73;
15'b0000100111110001101 : color = 12'he73;
15'b0000100111110001110 : color = 12'he73;
15'b0000100111110001111 : color = 12'he73;
15'b0000100111110010000 : color = 12'he73;
15'b0000100111110010001 : color = 12'he73;
15'b0000100111110010010 : color = 12'he73;
15'b0000100111110010011 : color = 12'he73;
15'b0000100111110010100 : color = 12'he73;
15'b0000100111110010101 : color = 12'he73;
15'b0000100111110010110 : color = 12'he73;
15'b0000100111110010111 : color = 12'he73;
15'b0000100111110011000 : color = 12'he73;
15'b0000100111110011001 : color = 12'he73;
15'b0000100111110011010 : color = 12'he73;
15'b0000100111110011011 : color = 12'he73;
15'b0000100111110011100 : color = 12'he73;
15'b0000100111110011101 : color = 12'he73;
15'b0000100111110011110 : color = 12'he73;
15'b0000100111110011111 : color = 12'he73;
15'b0000100111110100000 : color = 12'he73;
15'b0000100111110100001 : color = 12'he73;
15'b0000100111110100010 : color = 12'he73;
15'b0000100111110100011 : color = 12'he73;
15'b0000100111110100100 : color = 12'he73;
15'b0000100111110100101 : color = 12'he73;
15'b0000100111110100110 : color = 12'he73;
15'b0000100111110100111 : color = 12'he73;
15'b0000100111110101000 : color = 12'he73;
15'b0000100111110101001 : color = 12'he73;
15'b0000100111110101010 : color = 12'he73;
15'b0000100111110101011 : color = 12'he73;
15'b0000100111110101100 : color = 12'he73;
15'b0000100111110101101 : color = 12'he73;
15'b0000100111110101110 : color = 12'he73;
15'b0000100111110101111 : color = 12'he73;
15'b0000100111110110000 : color = 12'he73;
15'b0000100111110110001 : color = 12'he73;
15'b0000100111110110010 : color = 12'he73;
15'b0000100111110110011 : color = 12'he73;
15'b0000100111110110100 : color = 12'he73;
15'b0000100111110110101 : color = 12'he73;
15'b0000100111110110110 : color = 12'he73;
15'b0000100111110110111 : color = 12'he73;
15'b0000100111110111000 : color = 12'he73;
15'b0000100111110111001 : color = 12'he73;
15'b0000100111110111010 : color = 12'he73;
15'b0000100111110111011 : color = 12'he73;
15'b0000100111110111100 : color = 12'he73;
15'b0000100111110111101 : color = 12'he73;
15'b0000100111110111110 : color = 12'he73;
15'b0000100111110111111 : color = 12'he73;
15'b0000100111111000000 : color = 12'he73;
15'b0000100111111000001 : color = 12'he73;
15'b0000100111111000010 : color = 12'he73;
15'b0000100111111000011 : color = 12'he73;
15'b0000100111111000100 : color = 12'he73;
15'b0000100111111000101 : color = 12'he73;
15'b0000100111111000110 : color = 12'he73;
15'b0000100111111000111 : color = 12'he73;
15'b0000100111111001000 : color = 12'he73;
15'b0000100111111001001 : color = 12'he73;
15'b0000100111111001010 : color = 12'he73;
15'b0000100111111001011 : color = 12'he73;
15'b0000100111111001100 : color = 12'he73;
15'b0000100111111001101 : color = 12'he73;
15'b0000100111111001110 : color = 12'he73;
15'b0000100111111001111 : color = 12'he73;
15'b0000100111111010000 : color = 12'he73;
15'b0000100111111010001 : color = 12'he73;
15'b0000100111111010010 : color = 12'he73;
15'b0000100111111010011 : color = 12'he73;
15'b0000100111111010100 : color = 12'he73;
15'b0000100111111010101 : color = 12'he73;
15'b0000100111111010110 : color = 12'he73;
15'b0000100111111010111 : color = 12'he73;
15'b0000100111111011000 : color = 12'he73;
15'b0000100111111011001 : color = 12'he73;
15'b0000100111111011010 : color = 12'he73;
15'b0000100111111011011 : color = 12'he73;
15'b0000100111111011100 : color = 12'he73;
15'b0000100111111011101 : color = 12'he73;
15'b0000100111111011110 : color = 12'he73;
15'b0000100111111011111 : color = 12'he73;
15'b0000100111111100000 : color = 12'he73;
15'b0000100111111100001 : color = 12'he73;
15'b0000100111111100010 : color = 12'he73;
15'b0000100111111100011 : color = 12'he73;
15'b0000100111111100100 : color = 12'he73;
15'b0000100111111100101 : color = 12'he73;
15'b0000100111111100110 : color = 12'he73;
15'b0000100111111100111 : color = 12'he73;
15'b0000100111111101000 : color = 12'he73;
15'b0000100111111101001 : color = 12'he73;
15'b0000100111111101010 : color = 12'he73;
15'b0000100111111101011 : color = 12'he73;
15'b0000100111111101100 : color = 12'he73;
15'b0000100111111101101 : color = 12'he73;
15'b0000100111111101110 : color = 12'he73;
15'b0000100111111101111 : color = 12'he73;
15'b0000100111111110000 : color = 12'he73;
15'b0000100111111110001 : color = 12'he73;
15'b0000100111111110010 : color = 12'he73;
15'b0000100111111110011 : color = 12'he73;
15'b0000100111111110100 : color = 12'he73;
15'b0000100111111110101 : color = 12'he73;
15'b0000100111111110110 : color = 12'he73;
15'b0000100111111110111 : color = 12'he73;
15'b0000100111111111000 : color = 12'he73;
15'b0000100111111111001 : color = 12'he73;
15'b0000100111111111010 : color = 12'he73;
15'b0000100111111111011 : color = 12'he73;
15'b0000100111111111100 : color = 12'he73;
15'b0000100111111111101 : color = 12'he73;
15'b0000100111111111110 : color = 12'he73;
15'b0000100111111111111 : color = 12'he73;
15'b0000101000000000000 : color = 12'he73;
15'b0000101000000000001 : color = 12'he73;
15'b0000101000000000010 : color = 12'he73;
15'b0000101000000000011 : color = 12'he73;
15'b0000101000000000100 : color = 12'he73;
15'b0000101000000000101 : color = 12'he73;
15'b0000101000000000110 : color = 12'he73;
15'b0000101000000000111 : color = 12'he73;
15'b0000101000000001000 : color = 12'he73;
15'b0000101000000001001 : color = 12'he73;
15'b0000101000000001010 : color = 12'he73;
15'b0000101000000001011 : color = 12'he73;
15'b0000101000000001100 : color = 12'he73;
15'b0000101000000001101 : color = 12'he73;
15'b0000101000000001110 : color = 12'he73;
15'b0000101000000001111 : color = 12'he73;
15'b0000101000000010000 : color = 12'he73;
15'b0000101000000010001 : color = 12'he73;
15'b0000101000000010010 : color = 12'he73;
15'b0000101000000010011 : color = 12'he73;
15'b0000101000000010100 : color = 12'he73;
15'b0000101000000010101 : color = 12'he73;
15'b0000101000000010110 : color = 12'he73;
15'b0000101000000010111 : color = 12'he73;
15'b0000101000000011000 : color = 12'he73;
15'b0000101000000011001 : color = 12'he73;
15'b0000101000000011010 : color = 12'he73;
15'b0000101000000011011 : color = 12'he73;
15'b0000101000000011100 : color = 12'he73;
15'b0000101000000011101 : color = 12'he73;
15'b0000101000000011110 : color = 12'he73;
15'b0000101000000011111 : color = 12'he73;
15'b0000101000000100000 : color = 12'he73;
15'b0000101000000100001 : color = 12'he73;
15'b0000101000000100010 : color = 12'he73;
15'b0000101000000100011 : color = 12'he73;
15'b0000101000000100100 : color = 12'he73;
15'b0000101000000100101 : color = 12'he73;
15'b0000101000000100110 : color = 12'he73;
15'b0000101000000100111 : color = 12'he73;
15'b0000101000000101000 : color = 12'he73;
15'b0000101000000101001 : color = 12'he73;
15'b0000101000000101010 : color = 12'he73;
15'b0000101000000101011 : color = 12'he73;
15'b0000101000000101100 : color = 12'he73;
15'b0000101000000101101 : color = 12'he73;
15'b0000101000000101110 : color = 12'he73;
15'b0000101000000101111 : color = 12'he73;
15'b0000101000000110000 : color = 12'he73;
15'b0000101000000110001 : color = 12'he73;
15'b0000101000000110010 : color = 12'he73;
15'b0000101000000110011 : color = 12'he73;
15'b0000101000000110100 : color = 12'he73;
15'b0000101000000110101 : color = 12'he73;
15'b0000101000000110110 : color = 12'he73;
15'b0000101000000110111 : color = 12'he73;
15'b0000101000000111000 : color = 12'he73;
15'b0000101000000111001 : color = 12'he73;
15'b0000101000000111010 : color = 12'he73;
15'b0000101000000111011 : color = 12'he73;
15'b0000101000000111100 : color = 12'he73;
15'b0000101000000111101 : color = 12'he73;
15'b0000101000000111110 : color = 12'he73;
15'b0000101000000111111 : color = 12'he73;
15'b0000101000001000000 : color = 12'he73;
15'b0000101000001000001 : color = 12'he73;
15'b0000101000001000010 : color = 12'he73;
15'b0000101000001000011 : color = 12'he73;
15'b0000101000001000100 : color = 12'he73;
15'b0000101000001000101 : color = 12'he73;
15'b0000101000001000110 : color = 12'he73;
15'b0000101000001000111 : color = 12'he73;
15'b0000101000001001000 : color = 12'he73;
15'b0000101000001001001 : color = 12'he73;
15'b0000101000001001010 : color = 12'he73;
15'b0000101000001001011 : color = 12'he73;
15'b0000101000001001100 : color = 12'he73;
15'b0000101000001001101 : color = 12'he73;
15'b0000101000001001110 : color = 12'he73;
15'b0000101000001001111 : color = 12'he73;
15'b0000101000001010000 : color = 12'he73;
15'b0000101000001010001 : color = 12'he73;
15'b0000101000001010010 : color = 12'he73;
15'b0000101000001010011 : color = 12'he73;
15'b0000101000001010100 : color = 12'he73;
15'b0000101000001010101 : color = 12'he73;
15'b0000101000001010110 : color = 12'he73;
15'b0000101000001010111 : color = 12'he73;
15'b0000101000001011000 : color = 12'he73;
15'b0000101000001011001 : color = 12'he73;
15'b0000101000001011010 : color = 12'he73;
15'b0000101000001011011 : color = 12'he73;
15'b0000101000001011100 : color = 12'he73;
15'b0000101000001011101 : color = 12'he73;
15'b0000101000001011110 : color = 12'he73;
15'b0000101000001011111 : color = 12'he73;
15'b0000101000001100000 : color = 12'he73;
15'b0000101000001100001 : color = 12'he73;
15'b0000101000001100010 : color = 12'he73;
15'b0000101000001100011 : color = 12'he73;
15'b0000101000001100100 : color = 12'he73;
15'b0000101000001100101 : color = 12'he73;
15'b0000101000001100110 : color = 12'he73;
15'b0000101000001100111 : color = 12'he73;
15'b0000101000001101000 : color = 12'he73;
15'b0000101000001101001 : color = 12'he73;
15'b0000101000001101010 : color = 12'he73;
15'b0000101000001101011 : color = 12'he73;
15'b0000101000001101100 : color = 12'he73;
15'b0000101000001101101 : color = 12'he73;
15'b0000101000001101110 : color = 12'he73;
15'b0000101000001101111 : color = 12'he73;
15'b0000101000001110000 : color = 12'he73;
15'b0000101000001110001 : color = 12'he73;
15'b0000101000001110010 : color = 12'he73;
15'b0000101000001110011 : color = 12'he73;
15'b0000101000001110100 : color = 12'he73;
15'b0000101000001110101 : color = 12'he73;
15'b0000101000001110110 : color = 12'he73;
15'b0000101000001110111 : color = 12'he73;
15'b0000101000001111000 : color = 12'he73;
15'b0000101000001111001 : color = 12'he73;
15'b0000101000001111010 : color = 12'he73;
15'b0000101000001111011 : color = 12'he73;
15'b0000101000001111100 : color = 12'he73;
15'b0000101000001111101 : color = 12'he73;
15'b0000101000001111110 : color = 12'he73;
15'b0000101000001111111 : color = 12'he73;
15'b0000101000010000000 : color = 12'he73;
15'b0000101000010000001 : color = 12'he73;
15'b0000101000010000010 : color = 12'he73;
15'b0000101000010000011 : color = 12'he73;
15'b0000101000010000100 : color = 12'he73;
15'b0000101000010000101 : color = 12'he73;
15'b0000101000010000110 : color = 12'he73;
15'b0000101000010000111 : color = 12'he73;
15'b0000101000010001000 : color = 12'he73;
15'b0000101000010001001 : color = 12'he73;
15'b0000101000010001010 : color = 12'he73;
15'b0000101000010001011 : color = 12'he73;
15'b0000101000010001100 : color = 12'he73;
15'b0000101000010001101 : color = 12'he73;
15'b0000101000010001110 : color = 12'he73;
15'b0000101000010001111 : color = 12'he73;
15'b0000101000010010000 : color = 12'he73;
15'b0000101000010010001 : color = 12'he73;
15'b0000101000010010010 : color = 12'he73;
15'b0000101000010010011 : color = 12'he73;
15'b0000101000010010100 : color = 12'he73;
15'b0000101000010010101 : color = 12'he73;
15'b0000101000010010110 : color = 12'he73;
15'b0000101000010010111 : color = 12'he73;
15'b0000101000010011000 : color = 12'he73;
15'b0000101000010011001 : color = 12'he73;
15'b0000101000010011010 : color = 12'he73;
15'b0000101000010011011 : color = 12'he73;
15'b0000101000010011100 : color = 12'he73;
15'b0000101000010011101 : color = 12'he73;
15'b0000101000010011110 : color = 12'he73;
15'b0000101000010011111 : color = 12'he73;
15'b0000101000010100000 : color = 12'he73;
15'b0000101000010100001 : color = 12'he73;
15'b0000101000010100010 : color = 12'he73;
15'b0000101000010100011 : color = 12'he73;
15'b0000101000010100100 : color = 12'he73;
15'b0000101000010100101 : color = 12'he73;
15'b0000101000010100110 : color = 12'he73;
15'b0000101000010100111 : color = 12'he73;
15'b0000101000010101000 : color = 12'he73;
15'b0000101000010101001 : color = 12'he73;
15'b0000101000010101010 : color = 12'he73;
15'b0000101000010101011 : color = 12'he73;
15'b0000101000010101100 : color = 12'he73;
15'b0000101000010101101 : color = 12'he73;
15'b0000101000010101110 : color = 12'he73;
15'b0000101000010101111 : color = 12'he73;
15'b0000101000010110000 : color = 12'he73;
15'b0000101000010110001 : color = 12'he73;
15'b0000101000010110010 : color = 12'he73;
15'b0000101000010110011 : color = 12'he73;
15'b0000101000010110100 : color = 12'he73;
15'b0000101000010110101 : color = 12'he73;
15'b0000101000010110110 : color = 12'he73;
15'b0000101000010110111 : color = 12'he73;
15'b0000101000010111000 : color = 12'he73;
15'b0000101000010111001 : color = 12'he73;
15'b0000101000010111010 : color = 12'he73;
15'b0000101000010111011 : color = 12'he73;
15'b0000101000010111100 : color = 12'he73;
15'b0000101000010111101 : color = 12'he73;
15'b0000101000010111110 : color = 12'he73;
15'b0000101000010111111 : color = 12'he73;
15'b0000101000011000000 : color = 12'he73;
15'b0000101000011000001 : color = 12'he73;
15'b0000101000011000010 : color = 12'he73;
15'b0000101000011000011 : color = 12'he73;
15'b0000101000011000100 : color = 12'he73;
15'b0000101000011000101 : color = 12'he73;
15'b0000101000011000110 : color = 12'he73;
15'b0000101000011000111 : color = 12'he73;
15'b0000101000011001000 : color = 12'he73;
15'b0000101000011001001 : color = 12'he73;
15'b0000101000011001010 : color = 12'he73;
15'b0000101000011001011 : color = 12'he73;
15'b0000101000011001100 : color = 12'he73;
15'b0000101000011001101 : color = 12'he73;
15'b0000101000011001110 : color = 12'he73;
15'b0000101000011001111 : color = 12'he73;
15'b0000101000011010000 : color = 12'he73;
15'b0000101000011010001 : color = 12'he73;
15'b0000101000011010010 : color = 12'he73;
15'b0000101000011010011 : color = 12'he73;
15'b0000101000011010100 : color = 12'he73;
15'b0000101000011010101 : color = 12'he73;
15'b0000101000011010110 : color = 12'he73;
15'b0000101000011010111 : color = 12'he73;
15'b0000101000011011000 : color = 12'he73;
15'b0000101000011011001 : color = 12'he73;
15'b0000101000011011010 : color = 12'he73;
15'b0000101000011011011 : color = 12'he73;
15'b0000101000011011100 : color = 12'he73;
15'b0000101000011011101 : color = 12'he73;
15'b0000101000011011110 : color = 12'he73;
15'b0000101000011011111 : color = 12'he73;
15'b0000100111100011110 : color = 12'he73;
15'b0000100111100011111 : color = 12'he73;
15'b0000100111100100000 : color = 12'he73;
15'b0000100111100100001 : color = 12'he73;
15'b0000100111100100010 : color = 12'he73;
15'b0000100111100100011 : color = 12'he73;
15'b0000100111100100100 : color = 12'he73;
15'b0000100111100100101 : color = 12'he73;
15'b0000100111100100110 : color = 12'he73;
15'b0000100111100100111 : color = 12'he73;
15'b0000100111100101000 : color = 12'he73;
15'b0000100111100101001 : color = 12'he73;
15'b0000100111100101010 : color = 12'he73;
15'b0000100111100101011 : color = 12'he73;
15'b0000100111100101100 : color = 12'he73;
15'b0000100111100101101 : color = 12'he73;
15'b0000100111100101110 : color = 12'he73;
15'b0000100111100101111 : color = 12'he73;
15'b0000100111100110000 : color = 12'he73;
15'b0000100111100110001 : color = 12'he73;
15'b0000100111100110010 : color = 12'he73;
15'b0000100111100110011 : color = 12'he73;
15'b0000100111100110100 : color = 12'he73;
15'b0000100111100110101 : color = 12'he73;
15'b0000100111100110110 : color = 12'he73;
15'b0000100111100110111 : color = 12'he73;
15'b0000100111100111000 : color = 12'he73;
15'b0000100111100111001 : color = 12'he73;
15'b0000100111100111010 : color = 12'he73;
15'b0000100111100111011 : color = 12'he73;
15'b0000100111100111100 : color = 12'he73;
15'b0000100111100111101 : color = 12'he73;
15'b0000100111100111110 : color = 12'he73;
15'b0000100111100111111 : color = 12'he73;
15'b0000100111101000000 : color = 12'he73;
15'b0000100111101000001 : color = 12'he73;
15'b0000100111101000010 : color = 12'he73;
15'b0000100111101000011 : color = 12'he73;
15'b0000100111101000100 : color = 12'he73;
15'b0000100111101000101 : color = 12'he73;
15'b0000100111101000110 : color = 12'he73;
15'b0000100111101000111 : color = 12'he73;
15'b0000100111101001000 : color = 12'he73;
15'b0000100111101001001 : color = 12'he73;
15'b0000100111101001010 : color = 12'he73;
15'b0000100111101001011 : color = 12'he73;
15'b0000100111101001100 : color = 12'he73;
15'b0000100111101001101 : color = 12'he73;
15'b0000100111101001110 : color = 12'he73;
15'b0000100111101001111 : color = 12'he73;
15'b0000100111101010000 : color = 12'he73;
15'b0000100111101010001 : color = 12'he73;
15'b0000100111101010010 : color = 12'he73;
15'b0000100111101010011 : color = 12'he73;
15'b0000100111101010100 : color = 12'he73;
15'b0000100111101010101 : color = 12'he73;
15'b0000100111101010110 : color = 12'he73;
15'b0000100111101010111 : color = 12'he73;
15'b0000100111101011000 : color = 12'he73;
15'b0000100111101011001 : color = 12'he73;
15'b0000100111101011010 : color = 12'he73;
15'b0000100111101011011 : color = 12'he73;
15'b0000100111101011100 : color = 12'he73;
15'b0000100111101011101 : color = 12'he73;
15'b0000100111101011110 : color = 12'he73;
15'b0000100111101011111 : color = 12'he73;
15'b0000100111101100000 : color = 12'he73;
15'b0000100111101100001 : color = 12'he73;
15'b0000100111101100010 : color = 12'he73;
15'b0000100111101100011 : color = 12'he73;
15'b0000100111101100100 : color = 12'he73;
15'b0000100111101100101 : color = 12'he73;
15'b0000100111101100110 : color = 12'he73;
15'b0000100111101100111 : color = 12'he73;
15'b0000100111101101000 : color = 12'he73;
15'b0000100111101101001 : color = 12'he73;
15'b0000100111101101010 : color = 12'he73;
15'b0000100111101101011 : color = 12'he73;
15'b0000100111101101100 : color = 12'he73;
15'b0000100111101101101 : color = 12'he73;
15'b0000100111101101110 : color = 12'he73;
15'b0000100111101101111 : color = 12'he73;
15'b0000100111101110000 : color = 12'he73;
15'b0000100111101110001 : color = 12'he73;
15'b0000100111101110010 : color = 12'he73;
15'b0000100111101110011 : color = 12'he73;
15'b0000100111101110100 : color = 12'he73;
15'b0000100111101110101 : color = 12'he73;
15'b0000100111101110110 : color = 12'he73;
15'b0000100111101110111 : color = 12'he73;
15'b0000100111101111000 : color = 12'he73;
15'b0000100111101111001 : color = 12'he73;
15'b0000100111101111010 : color = 12'he73;
15'b0000100111101111011 : color = 12'he73;
15'b0000100111101111100 : color = 12'he73;
15'b0000100111101111101 : color = 12'he73;
15'b0000100111101111110 : color = 12'he73;
15'b0000100111101111111 : color = 12'he73;
15'b0000100111110000000 : color = 12'he73;
15'b0000100111110000001 : color = 12'he73;
15'b0000100111110000010 : color = 12'he73;
15'b0000100111110000011 : color = 12'he73;
15'b0000100111110000100 : color = 12'he73;
15'b0000100111110000101 : color = 12'he73;
15'b0000100111110000110 : color = 12'he73;
15'b0000100111110000111 : color = 12'he73;
15'b0000100111110001000 : color = 12'he73;
15'b0000100111110001001 : color = 12'he73;
15'b0000100111110001010 : color = 12'hf41;
15'b0000100111110001011 : color = 12'hf42;
15'b0000100111110001100 : color = 12'hf73;
15'b0000100111110001101 : color = 12'he73;
15'b0000100111110001110 : color = 12'he73;
15'b0000100111110001111 : color = 12'he73;
15'b0000100111110010000 : color = 12'he73;
15'b0000100111110010001 : color = 12'he73;
15'b0000100111110010010 : color = 12'he73;
15'b0000100111110010011 : color = 12'he73;
15'b0000100111110010100 : color = 12'he73;
15'b0000100111110010101 : color = 12'he73;
15'b0000100111110010110 : color = 12'he73;
15'b0000100111110010111 : color = 12'he73;
15'b0000100111110011000 : color = 12'he73;
15'b0000100111110011001 : color = 12'he73;
15'b0000100111110011010 : color = 12'he73;
15'b0000100111110011011 : color = 12'he73;
15'b0000100111110011100 : color = 12'he73;
15'b0000100111110011101 : color = 12'he73;
15'b0000100111110011110 : color = 12'he73;
15'b0000100111110011111 : color = 12'he73;
15'b0000100111110100000 : color = 12'he73;
15'b0000100111110100001 : color = 12'he73;
15'b0000100111110100010 : color = 12'he73;
15'b0000100111110100011 : color = 12'he73;
15'b0000100111110100100 : color = 12'he73;
15'b0000100111110100101 : color = 12'he73;
15'b0000100111110100110 : color = 12'he73;
15'b0000100111110100111 : color = 12'he73;
15'b0000100111110101000 : color = 12'he73;
15'b0000100111110101001 : color = 12'he73;
15'b0000100111110101010 : color = 12'he73;
15'b0000100111110101011 : color = 12'he73;
15'b0000100111110101100 : color = 12'he73;
15'b0000100111110101101 : color = 12'he73;
15'b0000100111110101110 : color = 12'he73;
15'b0000100111110101111 : color = 12'he73;
15'b0000100111110110000 : color = 12'he73;
15'b0000100111110110001 : color = 12'he73;
15'b0000100111110110010 : color = 12'he73;
15'b0000100111110110011 : color = 12'he73;
15'b0000100111110110100 : color = 12'he73;
15'b0000100111110110101 : color = 12'he73;
15'b0000100111110110110 : color = 12'he73;
15'b0000100111110110111 : color = 12'he73;
15'b0000100111110111000 : color = 12'he73;
15'b0000100111110111001 : color = 12'he73;
15'b0000100111110111010 : color = 12'he73;
15'b0000100111110111011 : color = 12'he73;
15'b0000100111110111100 : color = 12'he73;
15'b0000100111110111101 : color = 12'he73;
15'b0000100111110111110 : color = 12'he73;
15'b0000100111110111111 : color = 12'he73;
15'b0000100111111000000 : color = 12'he73;
15'b0000100111111000001 : color = 12'he73;
15'b0000100111111000010 : color = 12'he73;
15'b0000100111111000011 : color = 12'he73;
15'b0000100111111000100 : color = 12'he73;
15'b0000100111111000101 : color = 12'he73;
15'b0000100111111000110 : color = 12'he73;
15'b0000100111111000111 : color = 12'he73;
15'b0000100111111001000 : color = 12'he73;
15'b0000100111111001001 : color = 12'he73;
15'b0000100111111001010 : color = 12'he73;
15'b0000100111111001011 : color = 12'he73;
15'b0000100111111001100 : color = 12'he73;
15'b0000100111111001101 : color = 12'he73;
15'b0000100111111001110 : color = 12'he73;
15'b0000100111111001111 : color = 12'he73;
15'b0000100111111010000 : color = 12'he73;
15'b0000100111111010001 : color = 12'he73;
15'b0000100111111010010 : color = 12'he73;
15'b0000100111111010011 : color = 12'he73;
15'b0000100111111010100 : color = 12'he73;
15'b0000100111111010101 : color = 12'he73;
15'b0000100111111010110 : color = 12'he73;
15'b0000100111111010111 : color = 12'he73;
15'b0000100111111011000 : color = 12'he73;
15'b0000100111111011001 : color = 12'he73;
15'b0000100111111011010 : color = 12'he73;
15'b0000100111111011011 : color = 12'he73;
15'b0000100111111011100 : color = 12'he73;
15'b0000100111111011101 : color = 12'he73;
15'b0000100111111011110 : color = 12'he73;
15'b0000100111111011111 : color = 12'he73;
15'b0000100111111100000 : color = 12'he72;
15'b0000100111111100001 : color = 12'hf11;
15'b0000100111111100010 : color = 12'hf52;
15'b0000100111111100011 : color = 12'he73;
15'b0000100111111100100 : color = 12'he73;
15'b0000100111111100101 : color = 12'he73;
15'b0000100111111100110 : color = 12'he73;
15'b0000100111111100111 : color = 12'he73;
15'b0000100111111101000 : color = 12'he73;
15'b0000100111111101001 : color = 12'he73;
15'b0000100111111101010 : color = 12'he73;
15'b0000100111111101011 : color = 12'he73;
15'b0000100111111101100 : color = 12'he73;
15'b0000100111111101101 : color = 12'he73;
15'b0000100111111101110 : color = 12'he73;
15'b0000100111111101111 : color = 12'he73;
15'b0000100111111110000 : color = 12'he73;
15'b0000100111111110001 : color = 12'he73;
15'b0000100111111110010 : color = 12'he73;
15'b0000100111111110011 : color = 12'he73;
15'b0000100111111110100 : color = 12'he73;
15'b0000100111111110101 : color = 12'he73;
15'b0000100111111110110 : color = 12'he73;
15'b0000100111111110111 : color = 12'he73;
15'b0000100111111111000 : color = 12'he73;
15'b0000100111111111001 : color = 12'he73;
15'b0000100111111111010 : color = 12'he73;
15'b0000100111111111011 : color = 12'he73;
15'b0000100111111111100 : color = 12'he73;
15'b0000100111111111101 : color = 12'he73;
15'b0000100111111111110 : color = 12'he73;
15'b0000100111111111111 : color = 12'he73;
15'b0000101000000000000 : color = 12'he73;
15'b0000101000000000001 : color = 12'he73;
15'b0000101000000000010 : color = 12'he73;
15'b0000101000000000011 : color = 12'he73;
15'b0000101000000000100 : color = 12'he73;
15'b0000101000000000101 : color = 12'he73;
15'b0000101000000000110 : color = 12'he73;
15'b0000101000000000111 : color = 12'he73;
15'b0000101000000001000 : color = 12'he73;
15'b0000101000000001001 : color = 12'he73;
15'b0000101000000001010 : color = 12'he73;
15'b0000101000000001011 : color = 12'he73;
15'b0000101000000001100 : color = 12'he73;
15'b0000101000000001101 : color = 12'he73;
15'b0000101000000001110 : color = 12'he73;
15'b0000101000000001111 : color = 12'he73;
15'b0000101000000010000 : color = 12'he73;
15'b0000101000000010001 : color = 12'he73;
15'b0000101000000010010 : color = 12'he73;
15'b0000101000000010011 : color = 12'he73;
15'b0000101000000010100 : color = 12'he73;
15'b0000101000000010101 : color = 12'he73;
15'b0000101000000010110 : color = 12'he73;
15'b0000101000000010111 : color = 12'he73;
15'b0000101000000011000 : color = 12'he73;
15'b0000101000000011001 : color = 12'he73;
15'b0000101000000011010 : color = 12'he73;
15'b0000101000000011011 : color = 12'he73;
15'b0000101000000011100 : color = 12'he73;
15'b0000101000000011101 : color = 12'he73;
15'b0000101000000011110 : color = 12'he73;
15'b0000101000000011111 : color = 12'he73;
15'b0000101000000100000 : color = 12'he73;
15'b0000101000000100001 : color = 12'he73;
15'b0000101000000100010 : color = 12'he73;
15'b0000101000000100011 : color = 12'he73;
15'b0000101000000100100 : color = 12'he73;
15'b0000101000000100101 : color = 12'he73;
15'b0000101000000100110 : color = 12'he73;
15'b0000101000000100111 : color = 12'he73;
15'b0000101000000101000 : color = 12'he73;
15'b0000101000000101001 : color = 12'he73;
15'b0000101000000101010 : color = 12'he73;
15'b0000101000000101011 : color = 12'he73;
15'b0000101000000101100 : color = 12'he73;
15'b0000101000000101101 : color = 12'he73;
15'b0000101000000101110 : color = 12'he73;
15'b0000101000000101111 : color = 12'he73;
15'b0000101000000110000 : color = 12'he73;
15'b0000101000000110001 : color = 12'he73;
15'b0000101000000110010 : color = 12'he73;
15'b0000101000000110011 : color = 12'he73;
15'b0000101000000110100 : color = 12'he73;
15'b0000101000000110101 : color = 12'he73;
15'b0000101000000110110 : color = 12'he73;
15'b0000101000000110111 : color = 12'he73;
15'b0000101000000111000 : color = 12'he73;
15'b0000101000000111001 : color = 12'he73;
15'b0000101000000111010 : color = 12'he73;
15'b0000101000000111011 : color = 12'he73;
15'b0000101000000111100 : color = 12'he73;
15'b0000101000000111101 : color = 12'he73;
15'b0000101000000111110 : color = 12'he73;
15'b0000101000000111111 : color = 12'he73;
15'b0000101000001000000 : color = 12'he73;
15'b0000101000001000001 : color = 12'he73;
15'b0000101000001000010 : color = 12'he73;
15'b0000101000001000011 : color = 12'he73;
15'b0000101000001000100 : color = 12'he73;
15'b0000101000001000101 : color = 12'he73;
15'b0000101000001000110 : color = 12'he73;
15'b0000101000001000111 : color = 12'he73;
15'b0000101000001001000 : color = 12'he73;
15'b0000101000001001001 : color = 12'he73;
15'b0000101000001001010 : color = 12'he73;
15'b0000101000001001011 : color = 12'he73;
15'b0000101000001001100 : color = 12'he73;
15'b0000101000001001101 : color = 12'he73;
15'b0000101000001001110 : color = 12'he73;
15'b0000101000001001111 : color = 12'he73;
15'b0000101000001010000 : color = 12'he73;
15'b0000101000001010001 : color = 12'he73;
15'b0000101000001010010 : color = 12'he73;
15'b0000101000001010011 : color = 12'he73;
15'b0000101000001010100 : color = 12'he73;
15'b0000101000001010101 : color = 12'he73;
15'b0000101000001010110 : color = 12'he73;
15'b0000101000001010111 : color = 12'he73;
15'b0000101000001011000 : color = 12'he73;
15'b0000101000001011001 : color = 12'he73;
15'b0000101000001011010 : color = 12'he73;
15'b0000101000001011011 : color = 12'he73;
15'b0000101000001011100 : color = 12'he73;
15'b0000101000001011101 : color = 12'he73;
15'b0000101000001011110 : color = 12'he73;
15'b0000101000001011111 : color = 12'hf41;
15'b0000101000001100000 : color = 12'hf42;
15'b0000101000001100001 : color = 12'hf73;
15'b0000101000001100010 : color = 12'he73;
15'b0000101000001100011 : color = 12'he73;
15'b0000101000001100100 : color = 12'he73;
15'b0000101000001100101 : color = 12'he73;
15'b0000101000001100110 : color = 12'he73;
15'b0000101000001100111 : color = 12'he73;
15'b0000101000001101000 : color = 12'he73;
15'b0000101000001101001 : color = 12'he73;
15'b0000101000001101010 : color = 12'he51;
15'b0000101000001101011 : color = 12'hf52;
15'b0000101000001101100 : color = 12'he73;
15'b0000101000001101101 : color = 12'he73;
15'b0000101000001101110 : color = 12'he73;
15'b0000101000001101111 : color = 12'he73;
15'b0000101000001110000 : color = 12'he73;
15'b0000101000001110001 : color = 12'he73;
15'b0000101000001110010 : color = 12'he73;
15'b0000101000001110011 : color = 12'he73;
15'b0000101000001110100 : color = 12'he73;
15'b0000101000001110101 : color = 12'he73;
15'b0000101000001110110 : color = 12'he73;
15'b0000101000001110111 : color = 12'he73;
15'b0000101000001111000 : color = 12'he73;
15'b0000101000001111001 : color = 12'he73;
15'b0000101000001111010 : color = 12'he73;
15'b0000101000001111011 : color = 12'he73;
15'b0000101000001111100 : color = 12'he73;
15'b0000101000001111101 : color = 12'he73;
15'b0000101000001111110 : color = 12'he73;
15'b0000101000001111111 : color = 12'he73;
15'b0000101000010000000 : color = 12'he73;
15'b0000101000010000001 : color = 12'he73;
15'b0000101000010000010 : color = 12'he73;
15'b0000101000010000011 : color = 12'he73;
15'b0000101000010000100 : color = 12'he73;
15'b0000101000010000101 : color = 12'he73;
15'b0000101000010000110 : color = 12'he73;
15'b0000101000010000111 : color = 12'he73;
15'b0000101000010001000 : color = 12'he73;
15'b0000101000010001001 : color = 12'he73;
15'b0000101000010001010 : color = 12'he73;
15'b0000101000010001011 : color = 12'he73;
15'b0000101000010001100 : color = 12'he73;
15'b0000101000010001101 : color = 12'he73;
15'b0000101000010001110 : color = 12'he73;
15'b0000101000010001111 : color = 12'he73;
15'b0000101000010010000 : color = 12'he73;
15'b0000101000010010001 : color = 12'he73;
15'b0000101000010010010 : color = 12'he73;
15'b0000101000010010011 : color = 12'he73;
15'b0000101000010010100 : color = 12'he73;
15'b0000101000010010101 : color = 12'he73;
15'b0000101000010010110 : color = 12'he73;
15'b0000101000010010111 : color = 12'he73;
15'b0000101000010011000 : color = 12'he73;
15'b0000101000010011001 : color = 12'he73;
15'b0000101000010011010 : color = 12'he73;
15'b0000101000010011011 : color = 12'he73;
15'b0000101000010011100 : color = 12'he73;
15'b0000101000010011101 : color = 12'he73;
15'b0000101000010011110 : color = 12'he73;
15'b0000101000010011111 : color = 12'he73;
15'b0000101000010100000 : color = 12'he73;
15'b0000101000010100001 : color = 12'he73;
15'b0000101000010100010 : color = 12'he73;
15'b0000101000010100011 : color = 12'he73;
15'b0000101000010100100 : color = 12'he73;
15'b0000101000010100101 : color = 12'he73;
15'b0000101000010100110 : color = 12'he73;
15'b0000101000010100111 : color = 12'he73;
15'b0000101000010101000 : color = 12'he73;
15'b0000101000010101001 : color = 12'he73;
15'b0000101000010101010 : color = 12'he73;
15'b0000101000010101011 : color = 12'he73;
15'b0000101000010101100 : color = 12'he73;
15'b0000101000010101101 : color = 12'he73;
15'b0000101000010101110 : color = 12'he73;
15'b0000101000010101111 : color = 12'he73;
15'b0000101000010110000 : color = 12'he73;
15'b0000101000010110001 : color = 12'he73;
15'b0000101000010110010 : color = 12'he73;
15'b0000101000010110011 : color = 12'he73;
15'b0000101000010110100 : color = 12'he73;
15'b0000101000010110101 : color = 12'he73;
15'b0000101000010110110 : color = 12'he73;
15'b0000101000010110111 : color = 12'he73;
15'b0000101000010111000 : color = 12'he73;
15'b0000101000010111001 : color = 12'he73;
15'b0000101000010111010 : color = 12'he73;
15'b0000101000010111011 : color = 12'he73;
15'b0000101000010111100 : color = 12'he73;
15'b0000101000010111101 : color = 12'he73;
15'b0000101000010111110 : color = 12'he73;
15'b0000101000010111111 : color = 12'he73;
15'b0000101000011000000 : color = 12'he73;
15'b0000101000011000001 : color = 12'he73;
15'b0000101000011000010 : color = 12'he73;
15'b0000101000011000011 : color = 12'he73;
15'b0000101000011000100 : color = 12'he73;
15'b0000101000011000101 : color = 12'he72;
15'b0000101000011000110 : color = 12'hf41;
15'b0000101000011000111 : color = 12'hf10;
15'b0000101000011001000 : color = 12'hf53;
15'b0000101000011001001 : color = 12'he73;
15'b0000101000011001010 : color = 12'he73;
15'b0000101000011001011 : color = 12'he73;
15'b0000101000011001100 : color = 12'he73;
15'b0000101000011001101 : color = 12'he73;
15'b0000101000011001110 : color = 12'he73;
15'b0000101000011001111 : color = 12'he73;
15'b0000101000011010000 : color = 12'he73;
15'b0000101000011010001 : color = 12'he73;
15'b0000101000011010010 : color = 12'he73;
15'b0000101000011010011 : color = 12'he73;
15'b0000101000011010100 : color = 12'he73;
15'b0000101000011010101 : color = 12'he73;
15'b0000101000011010110 : color = 12'he73;
15'b0000101000011010111 : color = 12'he73;
15'b0000101000011011000 : color = 12'he73;
15'b0000101000011011001 : color = 12'he73;
15'b0000101000011011010 : color = 12'he73;
15'b0000101000011011011 : color = 12'he73;
15'b0000101000011011100 : color = 12'he73;
15'b0000101000011011101 : color = 12'he73;
15'b0000101000011011110 : color = 12'he73;
15'b0000101000011011111 : color = 12'he73;
15'b0000101000011100000 : color = 12'he73;
15'b0000101000011100001 : color = 12'he73;
15'b0000101000011100010 : color = 12'he73;
15'b0000101000011100011 : color = 12'he73;
15'b0000101000011100100 : color = 12'hf31;
15'b0000101000011100101 : color = 12'hf52;
15'b0000101000011100110 : color = 12'he73;
15'b0000101000011100111 : color = 12'he73;
15'b0000101000011101000 : color = 12'he73;
15'b0000101000011101001 : color = 12'he73;
15'b0000101000011101010 : color = 12'he73;
15'b0000101000011101011 : color = 12'he73;
15'b0000101000011101100 : color = 12'he73;
15'b0000101000011101101 : color = 12'he61;
15'b0000101000011101110 : color = 12'hf31;
15'b0000101000011101111 : color = 12'hf63;
15'b0000101000011110000 : color = 12'he73;
15'b0000101000011110001 : color = 12'he73;
15'b0000101000011110010 : color = 12'he73;
15'b0000101000011110011 : color = 12'he73;
15'b0000101000011110100 : color = 12'he73;
15'b0000101000011110101 : color = 12'he73;
15'b0000101000011110110 : color = 12'he73;
15'b0000101000011110111 : color = 12'he73;
15'b0000101000011111000 : color = 12'he73;
15'b0000101000011111001 : color = 12'he73;
15'b0000101000011111010 : color = 12'he73;
15'b0000101000011111011 : color = 12'he73;
15'b0000101000011111100 : color = 12'he73;
15'b0000101000011111101 : color = 12'he73;
15'b0000101000011111110 : color = 12'he73;
15'b0000101000011111111 : color = 12'he73;
15'b0000101000100000000 : color = 12'he73;
15'b0000101000100000001 : color = 12'he73;
15'b0000101000100000010 : color = 12'he73;
15'b0000101000100000011 : color = 12'he73;
15'b0000101000100000100 : color = 12'he73;
15'b0000101000100000101 : color = 12'he73;
15'b0000101000100000110 : color = 12'he73;
15'b0000101000100000111 : color = 12'he73;
15'b0000101000100001000 : color = 12'he73;
15'b0000100111101000111 : color = 12'he73;
15'b0000100111101001000 : color = 12'he73;
15'b0000100111101001001 : color = 12'he73;
15'b0000100111101001010 : color = 12'he73;
15'b0000100111101001011 : color = 12'he73;
15'b0000100111101001100 : color = 12'he73;
15'b0000100111101001101 : color = 12'he73;
15'b0000100111101001110 : color = 12'he73;
15'b0000100111101001111 : color = 12'he73;
15'b0000100111101010000 : color = 12'he73;
15'b0000100111101010001 : color = 12'he73;
15'b0000100111101010010 : color = 12'he73;
15'b0000100111101010011 : color = 12'he73;
15'b0000100111101010100 : color = 12'he73;
15'b0000100111101010101 : color = 12'he73;
15'b0000100111101010110 : color = 12'he73;
15'b0000100111101010111 : color = 12'he73;
15'b0000100111101011000 : color = 12'he73;
15'b0000100111101011001 : color = 12'he73;
15'b0000100111101011010 : color = 12'he73;
15'b0000100111101011011 : color = 12'he73;
15'b0000100111101011100 : color = 12'he73;
15'b0000100111101011101 : color = 12'he73;
15'b0000100111101011110 : color = 12'hf41;
15'b0000100111101011111 : color = 12'hf32;
15'b0000100111101100000 : color = 12'hf73;
15'b0000100111101100001 : color = 12'he73;
15'b0000100111101100010 : color = 12'he73;
15'b0000100111101100011 : color = 12'he73;
15'b0000100111101100100 : color = 12'he73;
15'b0000100111101100101 : color = 12'he73;
15'b0000100111101100110 : color = 12'he73;
15'b0000100111101100111 : color = 12'he73;
15'b0000100111101101000 : color = 12'he73;
15'b0000100111101101001 : color = 12'he73;
15'b0000100111101101010 : color = 12'he73;
15'b0000100111101101011 : color = 12'he73;
15'b0000100111101101100 : color = 12'he73;
15'b0000100111101101101 : color = 12'he73;
15'b0000100111101101110 : color = 12'he73;
15'b0000100111101101111 : color = 12'he73;
15'b0000100111101110000 : color = 12'he73;
15'b0000100111101110001 : color = 12'he73;
15'b0000100111101110010 : color = 12'he73;
15'b0000100111101110011 : color = 12'he73;
15'b0000100111101110100 : color = 12'he73;
15'b0000100111101110101 : color = 12'he73;
15'b0000100111101110110 : color = 12'he73;
15'b0000100111101110111 : color = 12'he73;
15'b0000100111101111000 : color = 12'he73;
15'b0000100111101111001 : color = 12'he73;
15'b0000100111101111010 : color = 12'he73;
15'b0000100111101111011 : color = 12'he73;
15'b0000100111101111100 : color = 12'he73;
15'b0000100111101111101 : color = 12'he73;
15'b0000100111101111110 : color = 12'he73;
15'b0000100111101111111 : color = 12'he73;
15'b0000100111110000000 : color = 12'he73;
15'b0000100111110000001 : color = 12'he73;
15'b0000100111110000010 : color = 12'he73;
15'b0000100111110000011 : color = 12'he73;
15'b0000100111110000100 : color = 12'he73;
15'b0000100111110000101 : color = 12'he73;
15'b0000100111110000110 : color = 12'he73;
15'b0000100111110000111 : color = 12'he73;
15'b0000100111110001000 : color = 12'he73;
15'b0000100111110001001 : color = 12'he73;
15'b0000100111110001010 : color = 12'he61;
15'b0000100111110001011 : color = 12'hf32;
15'b0000100111110001100 : color = 12'he73;
15'b0000100111110001101 : color = 12'he73;
15'b0000100111110001110 : color = 12'he73;
15'b0000100111110001111 : color = 12'he73;
15'b0000100111110010000 : color = 12'he73;
15'b0000100111110010001 : color = 12'he73;
15'b0000100111110010010 : color = 12'he73;
15'b0000100111110010011 : color = 12'he73;
15'b0000100111110010100 : color = 12'he73;
15'b0000100111110010101 : color = 12'he73;
15'b0000100111110010110 : color = 12'he73;
15'b0000100111110010111 : color = 12'he73;
15'b0000100111110011000 : color = 12'he73;
15'b0000100111110011001 : color = 12'he73;
15'b0000100111110011010 : color = 12'he73;
15'b0000100111110011011 : color = 12'he73;
15'b0000100111110011100 : color = 12'he73;
15'b0000100111110011101 : color = 12'he73;
15'b0000100111110011110 : color = 12'he73;
15'b0000100111110011111 : color = 12'he73;
15'b0000100111110100000 : color = 12'he73;
15'b0000100111110100001 : color = 12'he73;
15'b0000100111110100010 : color = 12'he73;
15'b0000100111110100011 : color = 12'he73;
15'b0000100111110100100 : color = 12'he73;
15'b0000100111110100101 : color = 12'he73;
15'b0000100111110100110 : color = 12'he73;
15'b0000100111110100111 : color = 12'he73;
15'b0000100111110101000 : color = 12'he73;
15'b0000100111110101001 : color = 12'he73;
15'b0000100111110101010 : color = 12'he73;
15'b0000100111110101011 : color = 12'he73;
15'b0000100111110101100 : color = 12'he73;
15'b0000100111110101101 : color = 12'he73;
15'b0000100111110101110 : color = 12'he73;
15'b0000100111110101111 : color = 12'he73;
15'b0000100111110110000 : color = 12'he73;
15'b0000100111110110001 : color = 12'he73;
15'b0000100111110110010 : color = 12'he73;
15'b0000100111110110011 : color = 12'hf40;
15'b0000100111110110100 : color = 12'hf00;
15'b0000100111110110101 : color = 12'hf01;
15'b0000100111110110110 : color = 12'hf63;
15'b0000100111110110111 : color = 12'he73;
15'b0000100111110111000 : color = 12'he73;
15'b0000100111110111001 : color = 12'he73;
15'b0000100111110111010 : color = 12'he73;
15'b0000100111110111011 : color = 12'he73;
15'b0000100111110111100 : color = 12'he73;
15'b0000100111110111101 : color = 12'he73;
15'b0000100111110111110 : color = 12'he73;
15'b0000100111110111111 : color = 12'he73;
15'b0000100111111000000 : color = 12'he73;
15'b0000100111111000001 : color = 12'he73;
15'b0000100111111000010 : color = 12'he73;
15'b0000100111111000011 : color = 12'he73;
15'b0000100111111000100 : color = 12'he73;
15'b0000100111111000101 : color = 12'he73;
15'b0000100111111000110 : color = 12'he73;
15'b0000100111111000111 : color = 12'he73;
15'b0000100111111001000 : color = 12'he73;
15'b0000100111111001001 : color = 12'he73;
15'b0000100111111001010 : color = 12'he73;
15'b0000100111111001011 : color = 12'he73;
15'b0000100111111001100 : color = 12'he73;
15'b0000100111111001101 : color = 12'he73;
15'b0000100111111001110 : color = 12'he73;
15'b0000100111111001111 : color = 12'he73;
15'b0000100111111010000 : color = 12'he73;
15'b0000100111111010001 : color = 12'he73;
15'b0000100111111010010 : color = 12'he73;
15'b0000100111111010011 : color = 12'he73;
15'b0000100111111010100 : color = 12'he73;
15'b0000100111111010101 : color = 12'he73;
15'b0000100111111010110 : color = 12'he73;
15'b0000100111111010111 : color = 12'he73;
15'b0000100111111011000 : color = 12'he73;
15'b0000100111111011001 : color = 12'he73;
15'b0000100111111011010 : color = 12'he73;
15'b0000100111111011011 : color = 12'he73;
15'b0000100111111011100 : color = 12'he73;
15'b0000100111111011101 : color = 12'he73;
15'b0000100111111011110 : color = 12'he73;
15'b0000100111111011111 : color = 12'he73;
15'b0000100111111100000 : color = 12'he73;
15'b0000100111111100001 : color = 12'he73;
15'b0000100111111100010 : color = 12'he73;
15'b0000100111111100011 : color = 12'he73;
15'b0000100111111100100 : color = 12'he73;
15'b0000100111111100101 : color = 12'he73;
15'b0000100111111100110 : color = 12'he73;
15'b0000100111111100111 : color = 12'he73;
15'b0000100111111101000 : color = 12'he73;
15'b0000100111111101001 : color = 12'he73;
15'b0000100111111101010 : color = 12'hf41;
15'b0000100111111101011 : color = 12'hf42;
15'b0000100111111101100 : color = 12'hf73;
15'b0000100111111101101 : color = 12'he73;
15'b0000100111111101110 : color = 12'he73;
15'b0000100111111101111 : color = 12'he73;
15'b0000100111111110000 : color = 12'he73;
15'b0000100111111110001 : color = 12'he73;
15'b0000100111111110010 : color = 12'he73;
15'b0000100111111110011 : color = 12'he73;
15'b0000100111111110100 : color = 12'he73;
15'b0000100111111110101 : color = 12'he73;
15'b0000100111111110110 : color = 12'he73;
15'b0000100111111110111 : color = 12'he73;
15'b0000100111111111000 : color = 12'he73;
15'b0000100111111111001 : color = 12'he73;
15'b0000100111111111010 : color = 12'he73;
15'b0000100111111111011 : color = 12'he73;
15'b0000100111111111100 : color = 12'he73;
15'b0000100111111111101 : color = 12'he73;
15'b0000100111111111110 : color = 12'he73;
15'b0000100111111111111 : color = 12'he73;
15'b0000101000000000000 : color = 12'he73;
15'b0000101000000000001 : color = 12'he73;
15'b0000101000000000010 : color = 12'he73;
15'b0000101000000000011 : color = 12'he73;
15'b0000101000000000100 : color = 12'he73;
15'b0000101000000000101 : color = 12'he73;
15'b0000101000000000110 : color = 12'he73;
15'b0000101000000000111 : color = 12'he73;
15'b0000101000000001000 : color = 12'he73;
15'b0000101000000001001 : color = 12'he73;
15'b0000101000000001010 : color = 12'he61;
15'b0000101000000001011 : color = 12'hf00;
15'b0000101000000001100 : color = 12'hf31;
15'b0000101000000001101 : color = 12'hf73;
15'b0000101000000001110 : color = 12'he73;
15'b0000101000000001111 : color = 12'he73;
15'b0000101000000010000 : color = 12'he73;
15'b0000101000000010001 : color = 12'he73;
15'b0000101000000010010 : color = 12'he73;
15'b0000101000000010011 : color = 12'he73;
15'b0000101000000010100 : color = 12'he73;
15'b0000101000000010101 : color = 12'he73;
15'b0000101000000010110 : color = 12'he73;
15'b0000101000000010111 : color = 12'he73;
15'b0000101000000011000 : color = 12'he73;
15'b0000101000000011001 : color = 12'he73;
15'b0000101000000011010 : color = 12'he73;
15'b0000101000000011011 : color = 12'he73;
15'b0000101000000011100 : color = 12'he73;
15'b0000101000000011101 : color = 12'he73;
15'b0000101000000011110 : color = 12'he73;
15'b0000101000000011111 : color = 12'he73;
15'b0000101000000100000 : color = 12'he73;
15'b0000101000000100001 : color = 12'he73;
15'b0000101000000100010 : color = 12'he73;
15'b0000101000000100011 : color = 12'he73;
15'b0000101000000100100 : color = 12'he73;
15'b0000101000000100101 : color = 12'he73;
15'b0000101000000100110 : color = 12'he73;
15'b0000101000000100111 : color = 12'he73;
15'b0000101000000101000 : color = 12'he73;
15'b0000101000000101001 : color = 12'he73;
15'b0000101000000101010 : color = 12'he73;
15'b0000101000000101011 : color = 12'he73;
15'b0000101000000101100 : color = 12'he73;
15'b0000101000000101101 : color = 12'he73;
15'b0000101000000101110 : color = 12'he73;
15'b0000101000000101111 : color = 12'he73;
15'b0000101000000110000 : color = 12'he73;
15'b0000101000000110001 : color = 12'he73;
15'b0000101000000110010 : color = 12'he73;
15'b0000101000000110011 : color = 12'he73;
15'b0000101000000110100 : color = 12'he73;
15'b0000101000000110101 : color = 12'he73;
15'b0000101000000110110 : color = 12'he73;
15'b0000101000000110111 : color = 12'he73;
15'b0000101000000111000 : color = 12'he73;
15'b0000101000000111001 : color = 12'he73;
15'b0000101000000111010 : color = 12'he73;
15'b0000101000000111011 : color = 12'he73;
15'b0000101000000111100 : color = 12'he73;
15'b0000101000000111101 : color = 12'he73;
15'b0000101000000111110 : color = 12'he73;
15'b0000101000000111111 : color = 12'he73;
15'b0000101000001000000 : color = 12'he51;
15'b0000101000001000001 : color = 12'hf42;
15'b0000101000001000010 : color = 12'he73;
15'b0000101000001000011 : color = 12'he73;
15'b0000101000001000100 : color = 12'he73;
15'b0000101000001000101 : color = 12'he73;
15'b0000101000001000110 : color = 12'he73;
15'b0000101000001000111 : color = 12'he73;
15'b0000101000001001000 : color = 12'he73;
15'b0000101000001001001 : color = 12'he73;
15'b0000101000001001010 : color = 12'he73;
15'b0000101000001001011 : color = 12'he73;
15'b0000101000001001100 : color = 12'he73;
15'b0000101000001001101 : color = 12'he73;
15'b0000101000001001110 : color = 12'he73;
15'b0000101000001001111 : color = 12'he73;
15'b0000101000001010000 : color = 12'he73;
15'b0000101000001010001 : color = 12'he73;
15'b0000101000001010010 : color = 12'he73;
15'b0000101000001010011 : color = 12'he73;
15'b0000101000001010100 : color = 12'he73;
15'b0000101000001010101 : color = 12'he73;
15'b0000101000001010110 : color = 12'he73;
15'b0000101000001010111 : color = 12'he73;
15'b0000101000001011000 : color = 12'he73;
15'b0000101000001011001 : color = 12'he73;
15'b0000101000001011010 : color = 12'he73;
15'b0000101000001011011 : color = 12'he73;
15'b0000101000001011100 : color = 12'hf30;
15'b0000101000001011101 : color = 12'hf42;
15'b0000101000001011110 : color = 12'hf73;
15'b0000101000001011111 : color = 12'he73;
15'b0000101000001100000 : color = 12'he73;
15'b0000101000001100001 : color = 12'he73;
15'b0000101000001100010 : color = 12'he73;
15'b0000101000001100011 : color = 12'he73;
15'b0000101000001100100 : color = 12'he73;
15'b0000101000001100101 : color = 12'he73;
15'b0000101000001100110 : color = 12'he73;
15'b0000101000001100111 : color = 12'he73;
15'b0000101000001101000 : color = 12'he73;
15'b0000101000001101001 : color = 12'he73;
15'b0000101000001101010 : color = 12'he73;
15'b0000101000001101011 : color = 12'he73;
15'b0000101000001101100 : color = 12'he73;
15'b0000101000001101101 : color = 12'he73;
15'b0000101000001101110 : color = 12'he73;
15'b0000101000001101111 : color = 12'he73;
15'b0000101000001110000 : color = 12'he73;
15'b0000101000001110001 : color = 12'he73;
15'b0000101000001110010 : color = 12'he73;
15'b0000101000001110011 : color = 12'he73;
15'b0000101000001110100 : color = 12'he73;
15'b0000101000001110101 : color = 12'he73;
15'b0000101000001110110 : color = 12'he73;
15'b0000101000001110111 : color = 12'he73;
15'b0000101000001111000 : color = 12'he73;
15'b0000101000001111001 : color = 12'he73;
15'b0000101000001111010 : color = 12'he73;
15'b0000101000001111011 : color = 12'he73;
15'b0000101000001111100 : color = 12'he73;
15'b0000101000001111101 : color = 12'he73;
15'b0000101000001111110 : color = 12'he73;
15'b0000101000001111111 : color = 12'he73;
15'b0000101000010000000 : color = 12'he73;
15'b0000101000010000001 : color = 12'he73;
15'b0000101000010000010 : color = 12'he73;
15'b0000101000010000011 : color = 12'he73;
15'b0000101000010000100 : color = 12'he73;
15'b0000101000010000101 : color = 12'he73;
15'b0000101000010000110 : color = 12'he73;
15'b0000101000010000111 : color = 12'he72;
15'b0000101000010001000 : color = 12'hf00;
15'b0000101000010001001 : color = 12'hf00;
15'b0000101000010001010 : color = 12'hf42;
15'b0000101000010001011 : color = 12'he73;
15'b0000101000010001100 : color = 12'he73;
15'b0000101000010001101 : color = 12'he73;
15'b0000101000010001110 : color = 12'he73;
15'b0000101000010001111 : color = 12'he73;
15'b0000101000010010000 : color = 12'he73;
15'b0000101000010010001 : color = 12'he73;
15'b0000101000010010010 : color = 12'he72;
15'b0000101000010010011 : color = 12'hf10;
15'b0000101000010010100 : color = 12'hf00;
15'b0000101000010010101 : color = 12'hf42;
15'b0000101000010010110 : color = 12'he73;
15'b0000101000010010111 : color = 12'he73;
15'b0000101000010011000 : color = 12'he73;
15'b0000101000010011001 : color = 12'he73;
15'b0000101000010011010 : color = 12'he73;
15'b0000101000010011011 : color = 12'he73;
15'b0000101000010011100 : color = 12'he73;
15'b0000101000010011101 : color = 12'he73;
15'b0000101000010011110 : color = 12'he73;
15'b0000101000010011111 : color = 12'he73;
15'b0000101000010100000 : color = 12'he73;
15'b0000101000010100001 : color = 12'he73;
15'b0000101000010100010 : color = 12'he73;
15'b0000101000010100011 : color = 12'he73;
15'b0000101000010100100 : color = 12'he73;
15'b0000101000010100101 : color = 12'he73;
15'b0000101000010100110 : color = 12'he73;
15'b0000101000010100111 : color = 12'he73;
15'b0000101000010101000 : color = 12'he73;
15'b0000101000010101001 : color = 12'he73;
15'b0000101000010101010 : color = 12'he73;
15'b0000101000010101011 : color = 12'he73;
15'b0000101000010101100 : color = 12'he73;
15'b0000101000010101101 : color = 12'he73;
15'b0000101000010101110 : color = 12'he73;
15'b0000101000010101111 : color = 12'he73;
15'b0000101000010110000 : color = 12'he73;
15'b0000101000010110001 : color = 12'he73;
15'b0000101000010110010 : color = 12'he73;
15'b0000101000010110011 : color = 12'he73;
15'b0000101000010110100 : color = 12'he73;
15'b0000101000010110101 : color = 12'he73;
15'b0000101000010110110 : color = 12'he73;
15'b0000101000010110111 : color = 12'he73;
15'b0000101000010111000 : color = 12'he73;
15'b0000101000010111001 : color = 12'he73;
15'b0000101000010111010 : color = 12'he73;
15'b0000101000010111011 : color = 12'he73;
15'b0000101000010111100 : color = 12'he73;
15'b0000101000010111101 : color = 12'he73;
15'b0000101000010111110 : color = 12'he73;
15'b0000101000010111111 : color = 12'he73;
15'b0000101000011000000 : color = 12'he73;
15'b0000101000011000001 : color = 12'he73;
15'b0000101000011000010 : color = 12'he73;
15'b0000101000011000011 : color = 12'he73;
15'b0000101000011000100 : color = 12'he73;
15'b0000101000011000101 : color = 12'he73;
15'b0000101000011000110 : color = 12'he73;
15'b0000101000011000111 : color = 12'he73;
15'b0000101000011001000 : color = 12'he73;
15'b0000101000011001001 : color = 12'he73;
15'b0000101000011001010 : color = 12'he73;
15'b0000101000011001011 : color = 12'he73;
15'b0000101000011001100 : color = 12'he73;
15'b0000101000011001101 : color = 12'he73;
15'b0000101000011001110 : color = 12'he73;
15'b0000101000011001111 : color = 12'he73;
15'b0000101000011010000 : color = 12'he73;
15'b0000101000011010001 : color = 12'he73;
15'b0000101000011010010 : color = 12'he73;
15'b0000101000011010011 : color = 12'he73;
15'b0000101000011010100 : color = 12'he73;
15'b0000101000011010101 : color = 12'he73;
15'b0000101000011010110 : color = 12'he73;
15'b0000101000011010111 : color = 12'he73;
15'b0000101000011011000 : color = 12'he73;
15'b0000101000011011001 : color = 12'he73;
15'b0000101000011011010 : color = 12'he73;
15'b0000101000011011011 : color = 12'he73;
15'b0000101000011011100 : color = 12'he73;
15'b0000101000011011101 : color = 12'he73;
15'b0000101000011011110 : color = 12'he73;
15'b0000101000011011111 : color = 12'he73;
15'b0000101000011100000 : color = 12'he73;
15'b0000101000011100001 : color = 12'he73;
15'b0000101000011100010 : color = 12'he73;
15'b0000101000011100011 : color = 12'he73;
15'b0000101000011100100 : color = 12'he73;
15'b0000101000011100101 : color = 12'he73;
15'b0000101000011100110 : color = 12'he73;
15'b0000101000011100111 : color = 12'he73;
15'b0000101000011101000 : color = 12'he73;
15'b0000101000011101001 : color = 12'he73;
15'b0000101000011101010 : color = 12'hf62;
15'b0000101000011101011 : color = 12'hf51;
15'b0000101000011101100 : color = 12'hf30;
15'b0000101000011101101 : color = 12'hf00;
15'b0000101000011101110 : color = 12'hf00;
15'b0000101000011101111 : color = 12'hf00;
15'b0000101000011110000 : color = 12'hf00;
15'b0000101000011110001 : color = 12'hf00;
15'b0000101000011110010 : color = 12'hf63;
15'b0000101000011110011 : color = 12'he73;
15'b0000101000011110100 : color = 12'he73;
15'b0000101000011110101 : color = 12'he73;
15'b0000101000011110110 : color = 12'he73;
15'b0000101000011110111 : color = 12'he73;
15'b0000101000011111000 : color = 12'he73;
15'b0000101000011111001 : color = 12'he73;
15'b0000101000011111010 : color = 12'he73;
15'b0000101000011111011 : color = 12'he73;
15'b0000101000011111100 : color = 12'he73;
15'b0000101000011111101 : color = 12'he73;
15'b0000101000011111110 : color = 12'he73;
15'b0000101000011111111 : color = 12'he73;
15'b0000101000100000000 : color = 12'he73;
15'b0000101000100000001 : color = 12'he73;
15'b0000101000100000010 : color = 12'he73;
15'b0000101000100000011 : color = 12'he73;
15'b0000101000100000100 : color = 12'he73;
15'b0000101000100000101 : color = 12'he73;
15'b0000101000100000110 : color = 12'he73;
15'b0000101000100000111 : color = 12'he73;
15'b0000101000100001000 : color = 12'he73;
15'b0000101000100001001 : color = 12'he73;
15'b0000101000100001010 : color = 12'he73;
15'b0000101000100001011 : color = 12'he73;
15'b0000101000100001100 : color = 12'he72;
15'b0000101000100001101 : color = 12'hf00;
15'b0000101000100001110 : color = 12'hf00;
15'b0000101000100001111 : color = 12'hf52;
15'b0000101000100010000 : color = 12'he73;
15'b0000101000100010001 : color = 12'he73;
15'b0000101000100010010 : color = 12'he73;
15'b0000101000100010011 : color = 12'he73;
15'b0000101000100010100 : color = 12'he73;
15'b0000101000100010101 : color = 12'he73;
15'b0000101000100010110 : color = 12'he73;
15'b0000101000100010111 : color = 12'hf40;
15'b0000101000100011000 : color = 12'hf00;
15'b0000101000100011001 : color = 12'hf42;
15'b0000101000100011010 : color = 12'he73;
15'b0000101000100011011 : color = 12'he73;
15'b0000101000100011100 : color = 12'he73;
15'b0000101000100011101 : color = 12'he73;
15'b0000101000100011110 : color = 12'he73;
15'b0000101000100011111 : color = 12'he73;
15'b0000101000100100000 : color = 12'he73;
15'b0000101000100100001 : color = 12'he73;
15'b0000101000100100010 : color = 12'he73;
15'b0000101000100100011 : color = 12'he73;
15'b0000101000100100100 : color = 12'he73;
15'b0000101000100100101 : color = 12'he73;
15'b0000101000100100110 : color = 12'he73;
15'b0000101000100100111 : color = 12'he73;
15'b0000101000100101000 : color = 12'he73;
15'b0000101000100101001 : color = 12'he73;
15'b0000101000100101010 : color = 12'he73;
15'b0000101000100101011 : color = 12'he73;
15'b0000101000100101100 : color = 12'he73;
15'b0000101000100101101 : color = 12'he73;
15'b0000101000100101110 : color = 12'he73;
15'b0000101000100101111 : color = 12'he73;
15'b0000101000100110000 : color = 12'he73;
15'b0000101000100110001 : color = 12'he73;
15'b0000100111101110000 : color = 12'he73;
15'b0000100111101110001 : color = 12'he73;
15'b0000100111101110010 : color = 12'he73;
15'b0000100111101110011 : color = 12'he73;
15'b0000100111101110100 : color = 12'he73;
15'b0000100111101110101 : color = 12'he73;
15'b0000100111101110110 : color = 12'he73;
15'b0000100111101110111 : color = 12'he73;
15'b0000100111101111000 : color = 12'he73;
15'b0000100111101111001 : color = 12'he73;
15'b0000100111101111010 : color = 12'he73;
15'b0000100111101111011 : color = 12'he73;
15'b0000100111101111100 : color = 12'he73;
15'b0000100111101111101 : color = 12'he73;
15'b0000100111101111110 : color = 12'he73;
15'b0000100111101111111 : color = 12'he73;
15'b0000100111110000000 : color = 12'he73;
15'b0000100111110000001 : color = 12'he73;
15'b0000100111110000010 : color = 12'he73;
15'b0000100111110000011 : color = 12'he73;
15'b0000100111110000100 : color = 12'he73;
15'b0000100111110000101 : color = 12'he73;
15'b0000100111110000110 : color = 12'he73;
15'b0000100111110000111 : color = 12'hf30;
15'b0000100111110001000 : color = 12'hf00;
15'b0000100111110001001 : color = 12'hf11;
15'b0000100111110001010 : color = 12'hf73;
15'b0000100111110001011 : color = 12'he73;
15'b0000100111110001100 : color = 12'he73;
15'b0000100111110001101 : color = 12'he73;
15'b0000100111110001110 : color = 12'he73;
15'b0000100111110001111 : color = 12'he73;
15'b0000100111110010000 : color = 12'he73;
15'b0000100111110010001 : color = 12'he73;
15'b0000100111110010010 : color = 12'he73;
15'b0000100111110010011 : color = 12'he73;
15'b0000100111110010100 : color = 12'he73;
15'b0000100111110010101 : color = 12'he73;
15'b0000100111110010110 : color = 12'he73;
15'b0000100111110010111 : color = 12'he73;
15'b0000100111110011000 : color = 12'he73;
15'b0000100111110011001 : color = 12'he73;
15'b0000100111110011010 : color = 12'he73;
15'b0000100111110011011 : color = 12'he73;
15'b0000100111110011100 : color = 12'he73;
15'b0000100111110011101 : color = 12'he73;
15'b0000100111110011110 : color = 12'he73;
15'b0000100111110011111 : color = 12'he73;
15'b0000100111110100000 : color = 12'he73;
15'b0000100111110100001 : color = 12'he73;
15'b0000100111110100010 : color = 12'he73;
15'b0000100111110100011 : color = 12'he73;
15'b0000100111110100100 : color = 12'he73;
15'b0000100111110100101 : color = 12'he73;
15'b0000100111110100110 : color = 12'he72;
15'b0000100111110100111 : color = 12'hf11;
15'b0000100111110101000 : color = 12'hf52;
15'b0000100111110101001 : color = 12'he73;
15'b0000100111110101010 : color = 12'he73;
15'b0000100111110101011 : color = 12'he73;
15'b0000100111110101100 : color = 12'he73;
15'b0000100111110101101 : color = 12'he73;
15'b0000100111110101110 : color = 12'he73;
15'b0000100111110101111 : color = 12'he73;
15'b0000100111110110000 : color = 12'he73;
15'b0000100111110110001 : color = 12'he73;
15'b0000100111110110010 : color = 12'hf41;
15'b0000100111110110011 : color = 12'hf00;
15'b0000100111110110100 : color = 12'hf00;
15'b0000100111110110101 : color = 12'hf42;
15'b0000100111110110110 : color = 12'he73;
15'b0000100111110110111 : color = 12'he73;
15'b0000100111110111000 : color = 12'he73;
15'b0000100111110111001 : color = 12'he73;
15'b0000100111110111010 : color = 12'he73;
15'b0000100111110111011 : color = 12'he73;
15'b0000100111110111100 : color = 12'he73;
15'b0000100111110111101 : color = 12'he73;
15'b0000100111110111110 : color = 12'he73;
15'b0000100111110111111 : color = 12'he73;
15'b0000100111111000000 : color = 12'he73;
15'b0000100111111000001 : color = 12'he73;
15'b0000100111111000010 : color = 12'he73;
15'b0000100111111000011 : color = 12'he73;
15'b0000100111111000100 : color = 12'he73;
15'b0000100111111000101 : color = 12'he73;
15'b0000100111111000110 : color = 12'he73;
15'b0000100111111000111 : color = 12'he73;
15'b0000100111111001000 : color = 12'he73;
15'b0000100111111001001 : color = 12'he73;
15'b0000100111111001010 : color = 12'he73;
15'b0000100111111001011 : color = 12'he73;
15'b0000100111111001100 : color = 12'he73;
15'b0000100111111001101 : color = 12'he73;
15'b0000100111111001110 : color = 12'he73;
15'b0000100111111001111 : color = 12'he73;
15'b0000100111111010000 : color = 12'he73;
15'b0000100111111010001 : color = 12'he73;
15'b0000100111111010010 : color = 12'he73;
15'b0000100111111010011 : color = 12'he73;
15'b0000100111111010100 : color = 12'he73;
15'b0000100111111010101 : color = 12'he73;
15'b0000100111111010110 : color = 12'he73;
15'b0000100111111010111 : color = 12'he73;
15'b0000100111111011000 : color = 12'he73;
15'b0000100111111011001 : color = 12'he73;
15'b0000100111111011010 : color = 12'he73;
15'b0000100111111011011 : color = 12'he73;
15'b0000100111111011100 : color = 12'hf40;
15'b0000100111111011101 : color = 12'hf00;
15'b0000100111111011110 : color = 12'hf53;
15'b0000100111111011111 : color = 12'he73;
15'b0000100111111100000 : color = 12'he73;
15'b0000100111111100001 : color = 12'he73;
15'b0000100111111100010 : color = 12'he73;
15'b0000100111111100011 : color = 12'he73;
15'b0000100111111100100 : color = 12'he73;
15'b0000100111111100101 : color = 12'he73;
15'b0000100111111100110 : color = 12'he73;
15'b0000100111111100111 : color = 12'he73;
15'b0000100111111101000 : color = 12'he73;
15'b0000100111111101001 : color = 12'he73;
15'b0000100111111101010 : color = 12'he73;
15'b0000100111111101011 : color = 12'he73;
15'b0000100111111101100 : color = 12'he73;
15'b0000100111111101101 : color = 12'he73;
15'b0000100111111101110 : color = 12'he73;
15'b0000100111111101111 : color = 12'he73;
15'b0000100111111110000 : color = 12'he73;
15'b0000100111111110001 : color = 12'he73;
15'b0000100111111110010 : color = 12'he73;
15'b0000100111111110011 : color = 12'he73;
15'b0000100111111110100 : color = 12'he73;
15'b0000100111111110101 : color = 12'he73;
15'b0000100111111110110 : color = 12'he73;
15'b0000100111111110111 : color = 12'he73;
15'b0000100111111111000 : color = 12'he73;
15'b0000100111111111001 : color = 12'he73;
15'b0000100111111111010 : color = 12'he73;
15'b0000100111111111011 : color = 12'he73;
15'b0000100111111111100 : color = 12'he73;
15'b0000100111111111101 : color = 12'he73;
15'b0000100111111111110 : color = 12'he73;
15'b0000100111111111111 : color = 12'he73;
15'b0000101000000000000 : color = 12'he73;
15'b0000101000000000001 : color = 12'he73;
15'b0000101000000000010 : color = 12'he73;
15'b0000101000000000011 : color = 12'he73;
15'b0000101000000000100 : color = 12'he73;
15'b0000101000000000101 : color = 12'he73;
15'b0000101000000000110 : color = 12'he73;
15'b0000101000000000111 : color = 12'he73;
15'b0000101000000001000 : color = 12'he73;
15'b0000101000000001001 : color = 12'he51;
15'b0000101000000001010 : color = 12'hf11;
15'b0000101000000001011 : color = 12'hf73;
15'b0000101000000001100 : color = 12'he73;
15'b0000101000000001101 : color = 12'he73;
15'b0000101000000001110 : color = 12'he73;
15'b0000101000000001111 : color = 12'he73;
15'b0000101000000010000 : color = 12'he73;
15'b0000101000000010001 : color = 12'he73;
15'b0000101000000010010 : color = 12'he73;
15'b0000101000000010011 : color = 12'hf40;
15'b0000101000000010100 : color = 12'hf00;
15'b0000101000000010101 : color = 12'hf42;
15'b0000101000000010110 : color = 12'he73;
15'b0000101000000010111 : color = 12'he73;
15'b0000101000000011000 : color = 12'he73;
15'b0000101000000011001 : color = 12'he73;
15'b0000101000000011010 : color = 12'he73;
15'b0000101000000011011 : color = 12'he73;
15'b0000101000000011100 : color = 12'he73;
15'b0000101000000011101 : color = 12'he73;
15'b0000101000000011110 : color = 12'he73;
15'b0000101000000011111 : color = 12'he73;
15'b0000101000000100000 : color = 12'he73;
15'b0000101000000100001 : color = 12'he73;
15'b0000101000000100010 : color = 12'he73;
15'b0000101000000100011 : color = 12'he73;
15'b0000101000000100100 : color = 12'he73;
15'b0000101000000100101 : color = 12'he73;
15'b0000101000000100110 : color = 12'he73;
15'b0000101000000100111 : color = 12'he73;
15'b0000101000000101000 : color = 12'he73;
15'b0000101000000101001 : color = 12'he73;
15'b0000101000000101010 : color = 12'he73;
15'b0000101000000101011 : color = 12'he73;
15'b0000101000000101100 : color = 12'he73;
15'b0000101000000101101 : color = 12'he73;
15'b0000101000000101110 : color = 12'he73;
15'b0000101000000101111 : color = 12'he73;
15'b0000101000000110000 : color = 12'he73;
15'b0000101000000110001 : color = 12'he73;
15'b0000101000000110010 : color = 12'he73;
15'b0000101000000110011 : color = 12'he73;
15'b0000101000000110100 : color = 12'hf40;
15'b0000101000000110101 : color = 12'hf00;
15'b0000101000000110110 : color = 12'hf11;
15'b0000101000000110111 : color = 12'hf73;
15'b0000101000000111000 : color = 12'he73;
15'b0000101000000111001 : color = 12'he73;
15'b0000101000000111010 : color = 12'he73;
15'b0000101000000111011 : color = 12'he73;
15'b0000101000000111100 : color = 12'he73;
15'b0000101000000111101 : color = 12'he73;
15'b0000101000000111110 : color = 12'he73;
15'b0000101000000111111 : color = 12'he73;
15'b0000101000001000000 : color = 12'he73;
15'b0000101000001000001 : color = 12'he73;
15'b0000101000001000010 : color = 12'he73;
15'b0000101000001000011 : color = 12'he73;
15'b0000101000001000100 : color = 12'he73;
15'b0000101000001000101 : color = 12'he73;
15'b0000101000001000110 : color = 12'he73;
15'b0000101000001000111 : color = 12'he73;
15'b0000101000001001000 : color = 12'he73;
15'b0000101000001001001 : color = 12'he73;
15'b0000101000001001010 : color = 12'he73;
15'b0000101000001001011 : color = 12'he73;
15'b0000101000001001100 : color = 12'he73;
15'b0000101000001001101 : color = 12'he73;
15'b0000101000001001110 : color = 12'he73;
15'b0000101000001001111 : color = 12'he73;
15'b0000101000001010000 : color = 12'he73;
15'b0000101000001010001 : color = 12'he73;
15'b0000101000001010010 : color = 12'he73;
15'b0000101000001010011 : color = 12'he73;
15'b0000101000001010100 : color = 12'he73;
15'b0000101000001010101 : color = 12'he73;
15'b0000101000001010110 : color = 12'hf41;
15'b0000101000001010111 : color = 12'hf42;
15'b0000101000001011000 : color = 12'hf73;
15'b0000101000001011001 : color = 12'he73;
15'b0000101000001011010 : color = 12'he73;
15'b0000101000001011011 : color = 12'he73;
15'b0000101000001011100 : color = 12'he73;
15'b0000101000001011101 : color = 12'he62;
15'b0000101000001011110 : color = 12'hf31;
15'b0000101000001011111 : color = 12'hf31;
15'b0000101000001100000 : color = 12'hf31;
15'b0000101000001100001 : color = 12'hf31;
15'b0000101000001100010 : color = 12'hf31;
15'b0000101000001100011 : color = 12'hf31;
15'b0000101000001100100 : color = 12'hf31;
15'b0000101000001100101 : color = 12'hf31;
15'b0000101000001100110 : color = 12'hf31;
15'b0000101000001100111 : color = 12'hf31;
15'b0000101000001101000 : color = 12'hf31;
15'b0000101000001101001 : color = 12'hf00;
15'b0000101000001101010 : color = 12'hf00;
15'b0000101000001101011 : color = 12'hf42;
15'b0000101000001101100 : color = 12'he73;
15'b0000101000001101101 : color = 12'he73;
15'b0000101000001101110 : color = 12'he73;
15'b0000101000001101111 : color = 12'he73;
15'b0000101000001110000 : color = 12'he73;
15'b0000101000001110001 : color = 12'he73;
15'b0000101000001110010 : color = 12'he73;
15'b0000101000001110011 : color = 12'he73;
15'b0000101000001110100 : color = 12'he73;
15'b0000101000001110101 : color = 12'he73;
15'b0000101000001110110 : color = 12'he73;
15'b0000101000001110111 : color = 12'he73;
15'b0000101000001111000 : color = 12'he73;
15'b0000101000001111001 : color = 12'he73;
15'b0000101000001111010 : color = 12'he73;
15'b0000101000001111011 : color = 12'he73;
15'b0000101000001111100 : color = 12'he73;
15'b0000101000001111101 : color = 12'he73;
15'b0000101000001111110 : color = 12'he73;
15'b0000101000001111111 : color = 12'he73;
15'b0000101000010000000 : color = 12'he73;
15'b0000101000010000001 : color = 12'he73;
15'b0000101000010000010 : color = 12'he73;
15'b0000101000010000011 : color = 12'he73;
15'b0000101000010000100 : color = 12'he73;
15'b0000101000010000101 : color = 12'hf30;
15'b0000101000010000110 : color = 12'hf00;
15'b0000101000010000111 : color = 12'hf52;
15'b0000101000010001000 : color = 12'he73;
15'b0000101000010001001 : color = 12'he73;
15'b0000101000010001010 : color = 12'he73;
15'b0000101000010001011 : color = 12'he73;
15'b0000101000010001100 : color = 12'he73;
15'b0000101000010001101 : color = 12'he73;
15'b0000101000010001110 : color = 12'he73;
15'b0000101000010001111 : color = 12'he73;
15'b0000101000010010000 : color = 12'he73;
15'b0000101000010010001 : color = 12'he73;
15'b0000101000010010010 : color = 12'he73;
15'b0000101000010010011 : color = 12'he73;
15'b0000101000010010100 : color = 12'he73;
15'b0000101000010010101 : color = 12'he73;
15'b0000101000010010110 : color = 12'he73;
15'b0000101000010010111 : color = 12'he73;
15'b0000101000010011000 : color = 12'he73;
15'b0000101000010011001 : color = 12'he73;
15'b0000101000010011010 : color = 12'he73;
15'b0000101000010011011 : color = 12'he73;
15'b0000101000010011100 : color = 12'he73;
15'b0000101000010011101 : color = 12'he73;
15'b0000101000010011110 : color = 12'he73;
15'b0000101000010011111 : color = 12'he73;
15'b0000101000010100000 : color = 12'he73;
15'b0000101000010100001 : color = 12'he73;
15'b0000101000010100010 : color = 12'he73;
15'b0000101000010100011 : color = 12'he73;
15'b0000101000010100100 : color = 12'he73;
15'b0000101000010100101 : color = 12'he73;
15'b0000101000010100110 : color = 12'he73;
15'b0000101000010100111 : color = 12'he73;
15'b0000101000010101000 : color = 12'he73;
15'b0000101000010101001 : color = 12'he73;
15'b0000101000010101010 : color = 12'he73;
15'b0000101000010101011 : color = 12'he73;
15'b0000101000010101100 : color = 12'he73;
15'b0000101000010101101 : color = 12'he73;
15'b0000101000010101110 : color = 12'he73;
15'b0000101000010101111 : color = 12'he73;
15'b0000101000010110000 : color = 12'hf40;
15'b0000101000010110001 : color = 12'hf00;
15'b0000101000010110010 : color = 12'hf53;
15'b0000101000010110011 : color = 12'he73;
15'b0000101000010110100 : color = 12'he73;
15'b0000101000010110101 : color = 12'he73;
15'b0000101000010110110 : color = 12'he73;
15'b0000101000010110111 : color = 12'he51;
15'b0000101000010111000 : color = 12'hf53;
15'b0000101000010111001 : color = 12'he73;
15'b0000101000010111010 : color = 12'he73;
15'b0000101000010111011 : color = 12'he51;
15'b0000101000010111100 : color = 12'hf00;
15'b0000101000010111101 : color = 12'hf53;
15'b0000101000010111110 : color = 12'he73;
15'b0000101000010111111 : color = 12'he73;
15'b0000101000011000000 : color = 12'he73;
15'b0000101000011000001 : color = 12'he73;
15'b0000101000011000010 : color = 12'he73;
15'b0000101000011000011 : color = 12'hf51;
15'b0000101000011000100 : color = 12'hf42;
15'b0000101000011000101 : color = 12'he73;
15'b0000101000011000110 : color = 12'he73;
15'b0000101000011000111 : color = 12'he73;
15'b0000101000011001000 : color = 12'he73;
15'b0000101000011001001 : color = 12'he73;
15'b0000101000011001010 : color = 12'he73;
15'b0000101000011001011 : color = 12'he73;
15'b0000101000011001100 : color = 12'he73;
15'b0000101000011001101 : color = 12'he73;
15'b0000101000011001110 : color = 12'he73;
15'b0000101000011001111 : color = 12'he73;
15'b0000101000011010000 : color = 12'he73;
15'b0000101000011010001 : color = 12'he73;
15'b0000101000011010010 : color = 12'he73;
15'b0000101000011010011 : color = 12'he73;
15'b0000101000011010100 : color = 12'he73;
15'b0000101000011010101 : color = 12'he73;
15'b0000101000011010110 : color = 12'he73;
15'b0000101000011010111 : color = 12'he73;
15'b0000101000011011000 : color = 12'he73;
15'b0000101000011011001 : color = 12'he73;
15'b0000101000011011010 : color = 12'he73;
15'b0000101000011011011 : color = 12'he73;
15'b0000101000011011100 : color = 12'he73;
15'b0000101000011011101 : color = 12'he73;
15'b0000101000011011110 : color = 12'he73;
15'b0000101000011011111 : color = 12'he73;
15'b0000101000011100000 : color = 12'he73;
15'b0000101000011100001 : color = 12'he73;
15'b0000101000011100010 : color = 12'he73;
15'b0000101000011100011 : color = 12'he51;
15'b0000101000011100100 : color = 12'hf63;
15'b0000101000011100101 : color = 12'he73;
15'b0000101000011100110 : color = 12'he73;
15'b0000101000011100111 : color = 12'he73;
15'b0000101000011101000 : color = 12'he73;
15'b0000101000011101001 : color = 12'he73;
15'b0000101000011101010 : color = 12'he73;
15'b0000101000011101011 : color = 12'he73;
15'b0000101000011101100 : color = 12'he73;
15'b0000101000011101101 : color = 12'he73;
15'b0000101000011101110 : color = 12'he72;
15'b0000101000011101111 : color = 12'hf11;
15'b0000101000011110000 : color = 12'hf63;
15'b0000101000011110001 : color = 12'he73;
15'b0000101000011110010 : color = 12'he73;
15'b0000101000011110011 : color = 12'he73;
15'b0000101000011110100 : color = 12'he73;
15'b0000101000011110101 : color = 12'he73;
15'b0000101000011110110 : color = 12'he73;
15'b0000101000011110111 : color = 12'he73;
15'b0000101000011111000 : color = 12'he73;
15'b0000101000011111001 : color = 12'he73;
15'b0000101000011111010 : color = 12'he73;
15'b0000101000011111011 : color = 12'he73;
15'b0000101000011111100 : color = 12'he73;
15'b0000101000011111101 : color = 12'he73;
15'b0000101000011111110 : color = 12'he73;
15'b0000101000011111111 : color = 12'he73;
15'b0000101000100000000 : color = 12'he73;
15'b0000101000100000001 : color = 12'he73;
15'b0000101000100000010 : color = 12'he73;
15'b0000101000100000011 : color = 12'he73;
15'b0000101000100000100 : color = 12'he73;
15'b0000101000100000101 : color = 12'he73;
15'b0000101000100000110 : color = 12'he73;
15'b0000101000100000111 : color = 12'he73;
15'b0000101000100001000 : color = 12'he73;
15'b0000101000100001001 : color = 12'he73;
15'b0000101000100001010 : color = 12'he73;
15'b0000101000100001011 : color = 12'he72;
15'b0000101000100001100 : color = 12'hf62;
15'b0000101000100001101 : color = 12'hf52;
15'b0000101000100001110 : color = 12'hf51;
15'b0000101000100001111 : color = 12'hf31;
15'b0000101000100010000 : color = 12'hf10;
15'b0000101000100010001 : color = 12'hf00;
15'b0000101000100010010 : color = 12'hf00;
15'b0000101000100010011 : color = 12'hf10;
15'b0000101000100010100 : color = 12'hf10;
15'b0000101000100010101 : color = 12'hf31;
15'b0000101000100010110 : color = 12'hf42;
15'b0000101000100010111 : color = 12'hf52;
15'b0000101000100011000 : color = 12'hf62;
15'b0000101000100011001 : color = 12'hf62;
15'b0000101000100011010 : color = 12'hf62;
15'b0000101000100011011 : color = 12'hf73;
15'b0000101000100011100 : color = 12'he73;
15'b0000101000100011101 : color = 12'he73;
15'b0000101000100011110 : color = 12'he73;
15'b0000101000100011111 : color = 12'he73;
15'b0000101000100100000 : color = 12'he73;
15'b0000101000100100001 : color = 12'he73;
15'b0000101000100100010 : color = 12'he73;
15'b0000101000100100011 : color = 12'he73;
15'b0000101000100100100 : color = 12'he73;
15'b0000101000100100101 : color = 12'he73;
15'b0000101000100100110 : color = 12'he73;
15'b0000101000100100111 : color = 12'he73;
15'b0000101000100101000 : color = 12'he73;
15'b0000101000100101001 : color = 12'he73;
15'b0000101000100101010 : color = 12'he73;
15'b0000101000100101011 : color = 12'he73;
15'b0000101000100101100 : color = 12'he73;
15'b0000101000100101101 : color = 12'he73;
15'b0000101000100101110 : color = 12'he73;
15'b0000101000100101111 : color = 12'he73;
15'b0000101000100110000 : color = 12'he73;
15'b0000101000100110001 : color = 12'he73;
15'b0000101000100110010 : color = 12'he73;
15'b0000101000100110011 : color = 12'he73;
15'b0000101000100110100 : color = 12'he73;
15'b0000101000100110101 : color = 12'hf40;
15'b0000101000100110110 : color = 12'hf00;
15'b0000101000100110111 : color = 12'hf42;
15'b0000101000100111000 : color = 12'he73;
15'b0000101000100111001 : color = 12'he73;
15'b0000101000100111010 : color = 12'he73;
15'b0000101000100111011 : color = 12'he73;
15'b0000101000100111100 : color = 12'he73;
15'b0000101000100111101 : color = 12'he73;
15'b0000101000100111110 : color = 12'he73;
15'b0000101000100111111 : color = 12'he73;
15'b0000101000101000000 : color = 12'he72;
15'b0000101000101000001 : color = 12'hf10;
15'b0000101000101000010 : color = 12'hf00;
15'b0000101000101000011 : color = 12'hf63;
15'b0000101000101000100 : color = 12'he73;
15'b0000101000101000101 : color = 12'he73;
15'b0000101000101000110 : color = 12'he73;
15'b0000101000101000111 : color = 12'he73;
15'b0000101000101001000 : color = 12'he73;
15'b0000101000101001001 : color = 12'he73;
15'b0000101000101001010 : color = 12'he73;
15'b0000101000101001011 : color = 12'he73;
15'b0000101000101001100 : color = 12'he73;
15'b0000101000101001101 : color = 12'he73;
15'b0000101000101001110 : color = 12'he73;
15'b0000101000101001111 : color = 12'he73;
15'b0000101000101010000 : color = 12'he73;
15'b0000101000101010001 : color = 12'he73;
15'b0000101000101010010 : color = 12'he73;
15'b0000101000101010011 : color = 12'he73;
15'b0000101000101010100 : color = 12'he73;
15'b0000101000101010101 : color = 12'he73;
15'b0000101000101010110 : color = 12'he73;
15'b0000101000101010111 : color = 12'he73;
15'b0000101000101011000 : color = 12'he73;
15'b0000101000101011001 : color = 12'he73;
15'b0000101000101011010 : color = 12'he73;
15'b0000100111110011001 : color = 12'he73;
15'b0000100111110011010 : color = 12'he73;
15'b0000100111110011011 : color = 12'he73;
15'b0000100111110011100 : color = 12'he73;
15'b0000100111110011101 : color = 12'he73;
15'b0000100111110011110 : color = 12'he73;
15'b0000100111110011111 : color = 12'he73;
15'b0000100111110100000 : color = 12'he73;
15'b0000100111110100001 : color = 12'he73;
15'b0000100111110100010 : color = 12'he73;
15'b0000100111110100011 : color = 12'he73;
15'b0000100111110100100 : color = 12'he73;
15'b0000100111110100101 : color = 12'he73;
15'b0000100111110100110 : color = 12'he73;
15'b0000100111110100111 : color = 12'he73;
15'b0000100111110101000 : color = 12'he73;
15'b0000100111110101001 : color = 12'he73;
15'b0000100111110101010 : color = 12'he51;
15'b0000100111110101011 : color = 12'hf31;
15'b0000100111110101100 : color = 12'hf73;
15'b0000100111110101101 : color = 12'he73;
15'b0000100111110101110 : color = 12'he73;
15'b0000100111110101111 : color = 12'he72;
15'b0000100111110110000 : color = 12'hf10;
15'b0000100111110110001 : color = 12'hf01;
15'b0000100111110110010 : color = 12'hf73;
15'b0000100111110110011 : color = 12'he73;
15'b0000100111110110100 : color = 12'he73;
15'b0000100111110110101 : color = 12'he73;
15'b0000100111110110110 : color = 12'he73;
15'b0000100111110110111 : color = 12'he73;
15'b0000100111110111000 : color = 12'he73;
15'b0000100111110111001 : color = 12'he73;
15'b0000100111110111010 : color = 12'he73;
15'b0000100111110111011 : color = 12'he73;
15'b0000100111110111100 : color = 12'he73;
15'b0000100111110111101 : color = 12'he73;
15'b0000100111110111110 : color = 12'he73;
15'b0000100111110111111 : color = 12'he73;
15'b0000100111111000000 : color = 12'he73;
15'b0000100111111000001 : color = 12'he73;
15'b0000100111111000010 : color = 12'he73;
15'b0000100111111000011 : color = 12'he73;
15'b0000100111111000100 : color = 12'he73;
15'b0000100111111000101 : color = 12'he73;
15'b0000100111111000110 : color = 12'he73;
15'b0000100111111000111 : color = 12'he73;
15'b0000100111111001000 : color = 12'he73;
15'b0000100111111001001 : color = 12'he73;
15'b0000100111111001010 : color = 12'he73;
15'b0000100111111001011 : color = 12'he73;
15'b0000100111111001100 : color = 12'he73;
15'b0000100111111001101 : color = 12'he73;
15'b0000100111111001110 : color = 12'he73;
15'b0000100111111001111 : color = 12'he73;
15'b0000100111111010000 : color = 12'he51;
15'b0000100111111010001 : color = 12'hf00;
15'b0000100111111010010 : color = 12'hf32;
15'b0000100111111010011 : color = 12'he73;
15'b0000100111111010100 : color = 12'he73;
15'b0000100111111010101 : color = 12'he73;
15'b0000100111111010110 : color = 12'he72;
15'b0000100111111010111 : color = 12'hf63;
15'b0000100111111011000 : color = 12'he73;
15'b0000100111111011001 : color = 12'hf51;
15'b0000100111111011010 : color = 12'hf10;
15'b0000100111111011011 : color = 12'hf11;
15'b0000100111111011100 : color = 12'hf52;
15'b0000100111111011101 : color = 12'hf73;
15'b0000100111111011110 : color = 12'he73;
15'b0000100111111011111 : color = 12'he73;
15'b0000100111111100000 : color = 12'he73;
15'b0000100111111100001 : color = 12'he73;
15'b0000100111111100010 : color = 12'he73;
15'b0000100111111100011 : color = 12'he73;
15'b0000100111111100100 : color = 12'he73;
15'b0000100111111100101 : color = 12'he73;
15'b0000100111111100110 : color = 12'he73;
15'b0000100111111100111 : color = 12'he73;
15'b0000100111111101000 : color = 12'he73;
15'b0000100111111101001 : color = 12'he73;
15'b0000100111111101010 : color = 12'he73;
15'b0000100111111101011 : color = 12'he73;
15'b0000100111111101100 : color = 12'he73;
15'b0000100111111101101 : color = 12'he73;
15'b0000100111111101110 : color = 12'he73;
15'b0000100111111101111 : color = 12'he73;
15'b0000100111111110000 : color = 12'he73;
15'b0000100111111110001 : color = 12'he73;
15'b0000100111111110010 : color = 12'he73;
15'b0000100111111110011 : color = 12'he73;
15'b0000100111111110100 : color = 12'he73;
15'b0000100111111110101 : color = 12'he73;
15'b0000100111111110110 : color = 12'he73;
15'b0000100111111110111 : color = 12'he73;
15'b0000100111111111000 : color = 12'he73;
15'b0000100111111111001 : color = 12'he73;
15'b0000100111111111010 : color = 12'he73;
15'b0000100111111111011 : color = 12'he73;
15'b0000100111111111100 : color = 12'he73;
15'b0000100111111111101 : color = 12'he73;
15'b0000100111111111110 : color = 12'he73;
15'b0000100111111111111 : color = 12'he73;
15'b0000101000000000000 : color = 12'he73;
15'b0000101000000000001 : color = 12'he73;
15'b0000101000000000010 : color = 12'he73;
15'b0000101000000000011 : color = 12'he73;
15'b0000101000000000100 : color = 12'he73;
15'b0000101000000000101 : color = 12'hf40;
15'b0000101000000000110 : color = 12'hf00;
15'b0000101000000000111 : color = 12'hf53;
15'b0000101000000001000 : color = 12'he73;
15'b0000101000000001001 : color = 12'he73;
15'b0000101000000001010 : color = 12'he73;
15'b0000101000000001011 : color = 12'he73;
15'b0000101000000001100 : color = 12'he73;
15'b0000101000000001101 : color = 12'he73;
15'b0000101000000001110 : color = 12'he73;
15'b0000101000000001111 : color = 12'he73;
15'b0000101000000010000 : color = 12'he73;
15'b0000101000000010001 : color = 12'he73;
15'b0000101000000010010 : color = 12'he73;
15'b0000101000000010011 : color = 12'he73;
15'b0000101000000010100 : color = 12'he73;
15'b0000101000000010101 : color = 12'he73;
15'b0000101000000010110 : color = 12'he73;
15'b0000101000000010111 : color = 12'he73;
15'b0000101000000011000 : color = 12'he73;
15'b0000101000000011001 : color = 12'he73;
15'b0000101000000011010 : color = 12'he73;
15'b0000101000000011011 : color = 12'he73;
15'b0000101000000011100 : color = 12'he73;
15'b0000101000000011101 : color = 12'he73;
15'b0000101000000011110 : color = 12'he73;
15'b0000101000000011111 : color = 12'he73;
15'b0000101000000100000 : color = 12'he73;
15'b0000101000000100001 : color = 12'he73;
15'b0000101000000100010 : color = 12'he73;
15'b0000101000000100011 : color = 12'he73;
15'b0000101000000100100 : color = 12'he73;
15'b0000101000000100101 : color = 12'he73;
15'b0000101000000100110 : color = 12'he62;
15'b0000101000000100111 : color = 12'hf31;
15'b0000101000000101000 : color = 12'hf31;
15'b0000101000000101001 : color = 12'hf31;
15'b0000101000000101010 : color = 12'hf31;
15'b0000101000000101011 : color = 12'hf31;
15'b0000101000000101100 : color = 12'hf31;
15'b0000101000000101101 : color = 12'hf31;
15'b0000101000000101110 : color = 12'hf31;
15'b0000101000000101111 : color = 12'hf31;
15'b0000101000000110000 : color = 12'hf31;
15'b0000101000000110001 : color = 12'hf30;
15'b0000101000000110010 : color = 12'hf00;
15'b0000101000000110011 : color = 12'hf00;
15'b0000101000000110100 : color = 12'hf11;
15'b0000101000000110101 : color = 12'hf73;
15'b0000101000000110110 : color = 12'he73;
15'b0000101000000110111 : color = 12'he73;
15'b0000101000000111000 : color = 12'he73;
15'b0000101000000111001 : color = 12'he73;
15'b0000101000000111010 : color = 12'he73;
15'b0000101000000111011 : color = 12'he73;
15'b0000101000000111100 : color = 12'hf40;
15'b0000101000000111101 : color = 12'hf01;
15'b0000101000000111110 : color = 12'hf73;
15'b0000101000000111111 : color = 12'he73;
15'b0000101000001000000 : color = 12'he73;
15'b0000101000001000001 : color = 12'he73;
15'b0000101000001000010 : color = 12'he73;
15'b0000101000001000011 : color = 12'he73;
15'b0000101000001000100 : color = 12'he73;
15'b0000101000001000101 : color = 12'he73;
15'b0000101000001000110 : color = 12'he73;
15'b0000101000001000111 : color = 12'he73;
15'b0000101000001001000 : color = 12'he73;
15'b0000101000001001001 : color = 12'he73;
15'b0000101000001001010 : color = 12'he73;
15'b0000101000001001011 : color = 12'he73;
15'b0000101000001001100 : color = 12'he73;
15'b0000101000001001101 : color = 12'he73;
15'b0000101000001001110 : color = 12'he73;
15'b0000101000001001111 : color = 12'he73;
15'b0000101000001010000 : color = 12'he73;
15'b0000101000001010001 : color = 12'he73;
15'b0000101000001010010 : color = 12'he73;
15'b0000101000001010011 : color = 12'he73;
15'b0000101000001010100 : color = 12'he73;
15'b0000101000001010101 : color = 12'he73;
15'b0000101000001010110 : color = 12'he73;
15'b0000101000001010111 : color = 12'he73;
15'b0000101000001011000 : color = 12'he73;
15'b0000101000001011001 : color = 12'he73;
15'b0000101000001011010 : color = 12'he73;
15'b0000101000001011011 : color = 12'he73;
15'b0000101000001011100 : color = 12'he73;
15'b0000101000001011101 : color = 12'he72;
15'b0000101000001011110 : color = 12'hf00;
15'b0000101000001011111 : color = 12'hf11;
15'b0000101000001100000 : color = 12'hf73;
15'b0000101000001100001 : color = 12'he73;
15'b0000101000001100010 : color = 12'he73;
15'b0000101000001100011 : color = 12'he73;
15'b0000101000001100100 : color = 12'he73;
15'b0000101000001100101 : color = 12'he73;
15'b0000101000001100110 : color = 12'he73;
15'b0000101000001100111 : color = 12'he73;
15'b0000101000001101000 : color = 12'he62;
15'b0000101000001101001 : color = 12'hf73;
15'b0000101000001101010 : color = 12'he73;
15'b0000101000001101011 : color = 12'he73;
15'b0000101000001101100 : color = 12'he73;
15'b0000101000001101101 : color = 12'he73;
15'b0000101000001101110 : color = 12'he73;
15'b0000101000001101111 : color = 12'he73;
15'b0000101000001110000 : color = 12'he73;
15'b0000101000001110001 : color = 12'he73;
15'b0000101000001110010 : color = 12'he73;
15'b0000101000001110011 : color = 12'he73;
15'b0000101000001110100 : color = 12'he73;
15'b0000101000001110101 : color = 12'he73;
15'b0000101000001110110 : color = 12'he73;
15'b0000101000001110111 : color = 12'he73;
15'b0000101000001111000 : color = 12'he73;
15'b0000101000001111001 : color = 12'he73;
15'b0000101000001111010 : color = 12'he73;
15'b0000101000001111011 : color = 12'he73;
15'b0000101000001111100 : color = 12'he73;
15'b0000101000001111101 : color = 12'he73;
15'b0000101000001111110 : color = 12'he73;
15'b0000101000001111111 : color = 12'he72;
15'b0000101000010000000 : color = 12'hf10;
15'b0000101000010000001 : color = 12'hf11;
15'b0000101000010000010 : color = 12'hf63;
15'b0000101000010000011 : color = 12'he73;
15'b0000101000010000100 : color = 12'he73;
15'b0000101000010000101 : color = 12'he73;
15'b0000101000010000110 : color = 12'he73;
15'b0000101000010000111 : color = 12'hf62;
15'b0000101000010001000 : color = 12'hf73;
15'b0000101000010001001 : color = 12'he73;
15'b0000101000010001010 : color = 12'he73;
15'b0000101000010001011 : color = 12'he73;
15'b0000101000010001100 : color = 12'he73;
15'b0000101000010001101 : color = 12'he73;
15'b0000101000010001110 : color = 12'he73;
15'b0000101000010001111 : color = 12'he73;
15'b0000101000010010000 : color = 12'he72;
15'b0000101000010010001 : color = 12'hf10;
15'b0000101000010010010 : color = 12'hf11;
15'b0000101000010010011 : color = 12'hf52;
15'b0000101000010010100 : color = 12'hf63;
15'b0000101000010010101 : color = 12'he73;
15'b0000101000010010110 : color = 12'he73;
15'b0000101000010010111 : color = 12'he73;
15'b0000101000010011000 : color = 12'he73;
15'b0000101000010011001 : color = 12'he73;
15'b0000101000010011010 : color = 12'he73;
15'b0000101000010011011 : color = 12'he73;
15'b0000101000010011100 : color = 12'he73;
15'b0000101000010011101 : color = 12'he73;
15'b0000101000010011110 : color = 12'he73;
15'b0000101000010011111 : color = 12'he73;
15'b0000101000010100000 : color = 12'he73;
15'b0000101000010100001 : color = 12'he73;
15'b0000101000010100010 : color = 12'he73;
15'b0000101000010100011 : color = 12'he73;
15'b0000101000010100100 : color = 12'he73;
15'b0000101000010100101 : color = 12'he73;
15'b0000101000010100110 : color = 12'he73;
15'b0000101000010100111 : color = 12'he73;
15'b0000101000010101000 : color = 12'he73;
15'b0000101000010101001 : color = 12'he73;
15'b0000101000010101010 : color = 12'he73;
15'b0000101000010101011 : color = 12'he73;
15'b0000101000010101100 : color = 12'he73;
15'b0000101000010101101 : color = 12'he73;
15'b0000101000010101110 : color = 12'hf30;
15'b0000101000010101111 : color = 12'hf01;
15'b0000101000010110000 : color = 12'hf73;
15'b0000101000010110001 : color = 12'he73;
15'b0000101000010110010 : color = 12'he73;
15'b0000101000010110011 : color = 12'he73;
15'b0000101000010110100 : color = 12'he73;
15'b0000101000010110101 : color = 12'he73;
15'b0000101000010110110 : color = 12'he73;
15'b0000101000010110111 : color = 12'he73;
15'b0000101000010111000 : color = 12'he73;
15'b0000101000010111001 : color = 12'he73;
15'b0000101000010111010 : color = 12'he73;
15'b0000101000010111011 : color = 12'he73;
15'b0000101000010111100 : color = 12'he73;
15'b0000101000010111101 : color = 12'he73;
15'b0000101000010111110 : color = 12'he73;
15'b0000101000010111111 : color = 12'he73;
15'b0000101000011000000 : color = 12'hf30;
15'b0000101000011000001 : color = 12'hf11;
15'b0000101000011000010 : color = 12'hf73;
15'b0000101000011000011 : color = 12'he73;
15'b0000101000011000100 : color = 12'he73;
15'b0000101000011000101 : color = 12'he73;
15'b0000101000011000110 : color = 12'he73;
15'b0000101000011000111 : color = 12'he73;
15'b0000101000011001000 : color = 12'he73;
15'b0000101000011001001 : color = 12'he73;
15'b0000101000011001010 : color = 12'he73;
15'b0000101000011001011 : color = 12'he73;
15'b0000101000011001100 : color = 12'he73;
15'b0000101000011001101 : color = 12'he73;
15'b0000101000011001110 : color = 12'he73;
15'b0000101000011001111 : color = 12'he73;
15'b0000101000011010000 : color = 12'he73;
15'b0000101000011010001 : color = 12'he73;
15'b0000101000011010010 : color = 12'he73;
15'b0000101000011010011 : color = 12'he73;
15'b0000101000011010100 : color = 12'he73;
15'b0000101000011010101 : color = 12'he73;
15'b0000101000011010110 : color = 12'he73;
15'b0000101000011010111 : color = 12'he73;
15'b0000101000011011000 : color = 12'he72;
15'b0000101000011011001 : color = 12'hf00;
15'b0000101000011011010 : color = 12'hf10;
15'b0000101000011011011 : color = 12'hf31;
15'b0000101000011011100 : color = 12'hf31;
15'b0000101000011011101 : color = 12'hf31;
15'b0000101000011011110 : color = 12'hf31;
15'b0000101000011011111 : color = 12'hf30;
15'b0000101000011100000 : color = 12'hf00;
15'b0000101000011100001 : color = 12'hf00;
15'b0000101000011100010 : color = 12'hf53;
15'b0000101000011100011 : color = 12'he72;
15'b0000101000011100100 : color = 12'hf10;
15'b0000101000011100101 : color = 12'hf10;
15'b0000101000011100110 : color = 12'hf31;
15'b0000101000011100111 : color = 12'hf31;
15'b0000101000011101000 : color = 12'hf31;
15'b0000101000011101001 : color = 12'hf31;
15'b0000101000011101010 : color = 12'hf31;
15'b0000101000011101011 : color = 12'hf30;
15'b0000101000011101100 : color = 12'hf00;
15'b0000101000011101101 : color = 12'hf00;
15'b0000101000011101110 : color = 12'hf52;
15'b0000101000011101111 : color = 12'he73;
15'b0000101000011110000 : color = 12'he73;
15'b0000101000011110001 : color = 12'he73;
15'b0000101000011110010 : color = 12'he73;
15'b0000101000011110011 : color = 12'he73;
15'b0000101000011110100 : color = 12'he73;
15'b0000101000011110101 : color = 12'he73;
15'b0000101000011110110 : color = 12'he73;
15'b0000101000011110111 : color = 12'he73;
15'b0000101000011111000 : color = 12'he73;
15'b0000101000011111001 : color = 12'he73;
15'b0000101000011111010 : color = 12'he73;
15'b0000101000011111011 : color = 12'he73;
15'b0000101000011111100 : color = 12'he73;
15'b0000101000011111101 : color = 12'he73;
15'b0000101000011111110 : color = 12'he73;
15'b0000101000011111111 : color = 12'he73;
15'b0000101000100000000 : color = 12'he73;
15'b0000101000100000001 : color = 12'he73;
15'b0000101000100000010 : color = 12'he73;
15'b0000101000100000011 : color = 12'he73;
15'b0000101000100000100 : color = 12'he73;
15'b0000101000100000101 : color = 12'he73;
15'b0000101000100000110 : color = 12'he73;
15'b0000101000100000111 : color = 12'he73;
15'b0000101000100001000 : color = 12'he73;
15'b0000101000100001001 : color = 12'hf40;
15'b0000101000100001010 : color = 12'hf32;
15'b0000101000100001011 : color = 12'he73;
15'b0000101000100001100 : color = 12'he51;
15'b0000101000100001101 : color = 12'hf00;
15'b0000101000100001110 : color = 12'hf31;
15'b0000101000100001111 : color = 12'hf31;
15'b0000101000100010000 : color = 12'hf31;
15'b0000101000100010001 : color = 12'hf31;
15'b0000101000100010010 : color = 12'hf31;
15'b0000101000100010011 : color = 12'hf31;
15'b0000101000100010100 : color = 12'hf31;
15'b0000101000100010101 : color = 12'hf31;
15'b0000101000100010110 : color = 12'hf31;
15'b0000101000100010111 : color = 12'hf10;
15'b0000101000100011000 : color = 12'hf00;
15'b0000101000100011001 : color = 12'hf32;
15'b0000101000100011010 : color = 12'hf73;
15'b0000101000100011011 : color = 12'he73;
15'b0000101000100011100 : color = 12'he73;
15'b0000101000100011101 : color = 12'he73;
15'b0000101000100011110 : color = 12'he73;
15'b0000101000100011111 : color = 12'he73;
15'b0000101000100100000 : color = 12'he73;
15'b0000101000100100001 : color = 12'he73;
15'b0000101000100100010 : color = 12'he73;
15'b0000101000100100011 : color = 12'he73;
15'b0000101000100100100 : color = 12'he73;
15'b0000101000100100101 : color = 12'he73;
15'b0000101000100100110 : color = 12'he73;
15'b0000101000100100111 : color = 12'he73;
15'b0000101000100101000 : color = 12'he73;
15'b0000101000100101001 : color = 12'he73;
15'b0000101000100101010 : color = 12'he73;
15'b0000101000100101011 : color = 12'he73;
15'b0000101000100101100 : color = 12'he73;
15'b0000101000100101101 : color = 12'he73;
15'b0000101000100101110 : color = 12'he73;
15'b0000101000100101111 : color = 12'he73;
15'b0000101000100110000 : color = 12'he51;
15'b0000101000100110001 : color = 12'hf41;
15'b0000101000100110010 : color = 12'hf31;
15'b0000101000100110011 : color = 12'hf31;
15'b0000101000100110100 : color = 12'hf31;
15'b0000101000100110101 : color = 12'hf31;
15'b0000101000100110110 : color = 12'hf52;
15'b0000101000100110111 : color = 12'hf52;
15'b0000101000100111000 : color = 12'hf52;
15'b0000101000100111001 : color = 12'hf51;
15'b0000101000100111010 : color = 12'hf11;
15'b0000101000100111011 : color = 12'hf52;
15'b0000101000100111100 : color = 12'he73;
15'b0000101000100111101 : color = 12'he73;
15'b0000101000100111110 : color = 12'he73;
15'b0000101000100111111 : color = 12'he73;
15'b0000101000101000000 : color = 12'he73;
15'b0000101000101000001 : color = 12'he73;
15'b0000101000101000010 : color = 12'he73;
15'b0000101000101000011 : color = 12'he73;
15'b0000101000101000100 : color = 12'he73;
15'b0000101000101000101 : color = 12'he73;
15'b0000101000101000110 : color = 12'he73;
15'b0000101000101000111 : color = 12'he73;
15'b0000101000101001000 : color = 12'he73;
15'b0000101000101001001 : color = 12'he73;
15'b0000101000101001010 : color = 12'he73;
15'b0000101000101001011 : color = 12'he73;
15'b0000101000101001100 : color = 12'he73;
15'b0000101000101001101 : color = 12'he73;
15'b0000101000101001110 : color = 12'he73;
15'b0000101000101001111 : color = 12'he73;
15'b0000101000101010000 : color = 12'he73;
15'b0000101000101010001 : color = 12'he73;
15'b0000101000101010010 : color = 12'he73;
15'b0000101000101010011 : color = 12'he73;
15'b0000101000101010100 : color = 12'he73;
15'b0000101000101010101 : color = 12'he73;
15'b0000101000101010110 : color = 12'he73;
15'b0000101000101010111 : color = 12'he73;
15'b0000101000101011000 : color = 12'he73;
15'b0000101000101011001 : color = 12'he73;
15'b0000101000101011010 : color = 12'he73;
15'b0000101000101011011 : color = 12'he73;
15'b0000101000101011100 : color = 12'he73;
15'b0000101000101011101 : color = 12'he72;
15'b0000101000101011110 : color = 12'hf10;
15'b0000101000101011111 : color = 12'hf11;
15'b0000101000101100000 : color = 12'hf73;
15'b0000101000101100001 : color = 12'he73;
15'b0000101000101100010 : color = 12'he73;
15'b0000101000101100011 : color = 12'he73;
15'b0000101000101100100 : color = 12'he73;
15'b0000101000101100101 : color = 12'he73;
15'b0000101000101100110 : color = 12'he73;
15'b0000101000101100111 : color = 12'he73;
15'b0000101000101101000 : color = 12'he73;
15'b0000101000101101001 : color = 12'he73;
15'b0000101000101101010 : color = 12'hf40;
15'b0000101000101101011 : color = 12'hf01;
15'b0000101000101101100 : color = 12'hf73;
15'b0000101000101101101 : color = 12'he73;
15'b0000101000101101110 : color = 12'he73;
15'b0000101000101101111 : color = 12'he73;
15'b0000101000101110000 : color = 12'hf40;
15'b0000101000101110001 : color = 12'hf11;
15'b0000101000101110010 : color = 12'hf73;
15'b0000101000101110011 : color = 12'he73;
15'b0000101000101110100 : color = 12'he73;
15'b0000101000101110101 : color = 12'he73;
15'b0000101000101110110 : color = 12'he73;
15'b0000101000101110111 : color = 12'he73;
15'b0000101000101111000 : color = 12'he73;
15'b0000101000101111001 : color = 12'he73;
15'b0000101000101111010 : color = 12'he73;
15'b0000101000101111011 : color = 12'he73;
15'b0000101000101111100 : color = 12'he73;
15'b0000101000101111101 : color = 12'he73;
15'b0000101000101111110 : color = 12'he73;
15'b0000101000101111111 : color = 12'he73;
15'b0000101000110000000 : color = 12'he73;
15'b0000101000110000001 : color = 12'he73;
15'b0000101000110000010 : color = 12'he73;
15'b0000101000110000011 : color = 12'he73;
15'b0000100111111000010 : color = 12'he73;
15'b0000100111111000011 : color = 12'he73;
15'b0000100111111000100 : color = 12'he73;
15'b0000100111111000101 : color = 12'he73;
15'b0000100111111000110 : color = 12'he73;
15'b0000100111111000111 : color = 12'he73;
15'b0000100111111001000 : color = 12'he73;
15'b0000100111111001001 : color = 12'he73;
15'b0000100111111001010 : color = 12'he61;
15'b0000100111111001011 : color = 12'hf31;
15'b0000100111111001100 : color = 12'hf31;
15'b0000100111111001101 : color = 12'hf31;
15'b0000100111111001110 : color = 12'hf31;
15'b0000100111111001111 : color = 12'hf31;
15'b0000100111111010000 : color = 12'hf31;
15'b0000100111111010001 : color = 12'hf31;
15'b0000100111111010010 : color = 12'hf31;
15'b0000100111111010011 : color = 12'hf00;
15'b0000100111111010100 : color = 12'hf00;
15'b0000100111111010101 : color = 12'hf32;
15'b0000100111111010110 : color = 12'hf73;
15'b0000100111111010111 : color = 12'he73;
15'b0000100111111011000 : color = 12'he72;
15'b0000100111111011001 : color = 12'hf00;
15'b0000100111111011010 : color = 12'hf32;
15'b0000100111111011011 : color = 12'he73;
15'b0000100111111011100 : color = 12'he73;
15'b0000100111111011101 : color = 12'he73;
15'b0000100111111011110 : color = 12'he73;
15'b0000100111111011111 : color = 12'he73;
15'b0000100111111100000 : color = 12'he73;
15'b0000100111111100001 : color = 12'he73;
15'b0000100111111100010 : color = 12'he73;
15'b0000100111111100011 : color = 12'he73;
15'b0000100111111100100 : color = 12'he73;
15'b0000100111111100101 : color = 12'he73;
15'b0000100111111100110 : color = 12'he73;
15'b0000100111111100111 : color = 12'he73;
15'b0000100111111101000 : color = 12'he73;
15'b0000100111111101001 : color = 12'he73;
15'b0000100111111101010 : color = 12'he73;
15'b0000100111111101011 : color = 12'he73;
15'b0000100111111101100 : color = 12'he73;
15'b0000100111111101101 : color = 12'he73;
15'b0000100111111101110 : color = 12'he73;
15'b0000100111111101111 : color = 12'he73;
15'b0000100111111110000 : color = 12'he73;
15'b0000100111111110001 : color = 12'he73;
15'b0000100111111110010 : color = 12'he73;
15'b0000100111111110011 : color = 12'he73;
15'b0000100111111110100 : color = 12'he73;
15'b0000100111111110101 : color = 12'he73;
15'b0000100111111110110 : color = 12'he73;
15'b0000100111111110111 : color = 12'he73;
15'b0000100111111111000 : color = 12'he73;
15'b0000100111111111001 : color = 12'he73;
15'b0000100111111111010 : color = 12'hf30;
15'b0000100111111111011 : color = 12'hf00;
15'b0000100111111111100 : color = 12'hf42;
15'b0000100111111111101 : color = 12'he73;
15'b0000100111111111110 : color = 12'he73;
15'b0000100111111111111 : color = 12'he61;
15'b0000101000000000000 : color = 12'hf00;
15'b0000101000000000001 : color = 12'hf11;
15'b0000101000000000010 : color = 12'hf52;
15'b0000101000000000011 : color = 12'hf73;
15'b0000101000000000100 : color = 12'he73;
15'b0000101000000000101 : color = 12'he73;
15'b0000101000000000110 : color = 12'he72;
15'b0000101000000000111 : color = 12'hf52;
15'b0000101000000001000 : color = 12'he73;
15'b0000101000000001001 : color = 12'he73;
15'b0000101000000001010 : color = 12'he73;
15'b0000101000000001011 : color = 12'he73;
15'b0000101000000001100 : color = 12'he73;
15'b0000101000000001101 : color = 12'he51;
15'b0000101000000001110 : color = 12'hf63;
15'b0000101000000001111 : color = 12'he73;
15'b0000101000000010000 : color = 12'he73;
15'b0000101000000010001 : color = 12'he73;
15'b0000101000000010010 : color = 12'he73;
15'b0000101000000010011 : color = 12'he73;
15'b0000101000000010100 : color = 12'he73;
15'b0000101000000010101 : color = 12'he73;
15'b0000101000000010110 : color = 12'he73;
15'b0000101000000010111 : color = 12'he73;
15'b0000101000000011000 : color = 12'he73;
15'b0000101000000011001 : color = 12'he73;
15'b0000101000000011010 : color = 12'he73;
15'b0000101000000011011 : color = 12'he73;
15'b0000101000000011100 : color = 12'he73;
15'b0000101000000011101 : color = 12'he73;
15'b0000101000000011110 : color = 12'he73;
15'b0000101000000011111 : color = 12'he73;
15'b0000101000000100000 : color = 12'he73;
15'b0000101000000100001 : color = 12'he73;
15'b0000101000000100010 : color = 12'he73;
15'b0000101000000100011 : color = 12'he73;
15'b0000101000000100100 : color = 12'he73;
15'b0000101000000100101 : color = 12'he73;
15'b0000101000000100110 : color = 12'he73;
15'b0000101000000100111 : color = 12'he73;
15'b0000101000000101000 : color = 12'he73;
15'b0000101000000101001 : color = 12'he73;
15'b0000101000000101010 : color = 12'he73;
15'b0000101000000101011 : color = 12'he73;
15'b0000101000000101100 : color = 12'he73;
15'b0000101000000101101 : color = 12'he73;
15'b0000101000000101110 : color = 12'he51;
15'b0000101000000101111 : color = 12'hf00;
15'b0000101000000110000 : color = 12'hf53;
15'b0000101000000110001 : color = 12'he73;
15'b0000101000000110010 : color = 12'he73;
15'b0000101000000110011 : color = 12'he73;
15'b0000101000000110100 : color = 12'he73;
15'b0000101000000110101 : color = 12'he73;
15'b0000101000000110110 : color = 12'he73;
15'b0000101000000110111 : color = 12'he72;
15'b0000101000000111000 : color = 12'hf10;
15'b0000101000000111001 : color = 12'hf42;
15'b0000101000000111010 : color = 12'he73;
15'b0000101000000111011 : color = 12'he73;
15'b0000101000000111100 : color = 12'he73;
15'b0000101000000111101 : color = 12'he73;
15'b0000101000000111110 : color = 12'he73;
15'b0000101000000111111 : color = 12'he73;
15'b0000101000001000000 : color = 12'he73;
15'b0000101000001000001 : color = 12'he73;
15'b0000101000001000010 : color = 12'he73;
15'b0000101000001000011 : color = 12'he73;
15'b0000101000001000100 : color = 12'he73;
15'b0000101000001000101 : color = 12'he73;
15'b0000101000001000110 : color = 12'he73;
15'b0000101000001000111 : color = 12'he73;
15'b0000101000001001000 : color = 12'he73;
15'b0000101000001001001 : color = 12'he73;
15'b0000101000001001010 : color = 12'he73;
15'b0000101000001001011 : color = 12'he73;
15'b0000101000001001100 : color = 12'he73;
15'b0000101000001001101 : color = 12'he73;
15'b0000101000001001110 : color = 12'he73;
15'b0000101000001001111 : color = 12'he73;
15'b0000101000001010000 : color = 12'hf62;
15'b0000101000001010001 : color = 12'hf73;
15'b0000101000001010010 : color = 12'he73;
15'b0000101000001010011 : color = 12'he73;
15'b0000101000001010100 : color = 12'he73;
15'b0000101000001010101 : color = 12'he61;
15'b0000101000001010110 : color = 12'hf00;
15'b0000101000001010111 : color = 12'hf52;
15'b0000101000001011000 : color = 12'he73;
15'b0000101000001011001 : color = 12'he73;
15'b0000101000001011010 : color = 12'he73;
15'b0000101000001011011 : color = 12'he73;
15'b0000101000001011100 : color = 12'he73;
15'b0000101000001011101 : color = 12'he73;
15'b0000101000001011110 : color = 12'he73;
15'b0000101000001011111 : color = 12'he73;
15'b0000101000001100000 : color = 12'he73;
15'b0000101000001100001 : color = 12'he73;
15'b0000101000001100010 : color = 12'he73;
15'b0000101000001100011 : color = 12'he73;
15'b0000101000001100100 : color = 12'he73;
15'b0000101000001100101 : color = 12'hf40;
15'b0000101000001100110 : color = 12'hf01;
15'b0000101000001100111 : color = 12'hf73;
15'b0000101000001101000 : color = 12'he73;
15'b0000101000001101001 : color = 12'he73;
15'b0000101000001101010 : color = 12'he73;
15'b0000101000001101011 : color = 12'he73;
15'b0000101000001101100 : color = 12'he73;
15'b0000101000001101101 : color = 12'he73;
15'b0000101000001101110 : color = 12'he73;
15'b0000101000001101111 : color = 12'he73;
15'b0000101000001110000 : color = 12'he73;
15'b0000101000001110001 : color = 12'he73;
15'b0000101000001110010 : color = 12'he73;
15'b0000101000001110011 : color = 12'he73;
15'b0000101000001110100 : color = 12'he73;
15'b0000101000001110101 : color = 12'he73;
15'b0000101000001110110 : color = 12'he73;
15'b0000101000001110111 : color = 12'he73;
15'b0000101000001111000 : color = 12'he73;
15'b0000101000001111001 : color = 12'he73;
15'b0000101000001111010 : color = 12'he73;
15'b0000101000001111011 : color = 12'he73;
15'b0000101000001111100 : color = 12'he73;
15'b0000101000001111101 : color = 12'he73;
15'b0000101000001111110 : color = 12'he73;
15'b0000101000001111111 : color = 12'he73;
15'b0000101000010000000 : color = 12'he73;
15'b0000101000010000001 : color = 12'he73;
15'b0000101000010000010 : color = 12'he73;
15'b0000101000010000011 : color = 12'he73;
15'b0000101000010000100 : color = 12'he73;
15'b0000101000010000101 : color = 12'he73;
15'b0000101000010000110 : color = 12'he73;
15'b0000101000010000111 : color = 12'hf41;
15'b0000101000010001000 : color = 12'hf63;
15'b0000101000010001001 : color = 12'he73;
15'b0000101000010001010 : color = 12'he73;
15'b0000101000010001011 : color = 12'he73;
15'b0000101000010001100 : color = 12'he73;
15'b0000101000010001101 : color = 12'he73;
15'b0000101000010001110 : color = 12'he73;
15'b0000101000010001111 : color = 12'he73;
15'b0000101000010010000 : color = 12'he61;
15'b0000101000010010001 : color = 12'hf00;
15'b0000101000010010010 : color = 12'hf11;
15'b0000101000010010011 : color = 12'hf73;
15'b0000101000010010100 : color = 12'he73;
15'b0000101000010010101 : color = 12'he73;
15'b0000101000010010110 : color = 12'he73;
15'b0000101000010010111 : color = 12'he73;
15'b0000101000010011000 : color = 12'he73;
15'b0000101000010011001 : color = 12'he73;
15'b0000101000010011010 : color = 12'he73;
15'b0000101000010011011 : color = 12'he73;
15'b0000101000010011100 : color = 12'he73;
15'b0000101000010011101 : color = 12'he73;
15'b0000101000010011110 : color = 12'he73;
15'b0000101000010011111 : color = 12'he73;
15'b0000101000010100000 : color = 12'he73;
15'b0000101000010100001 : color = 12'he73;
15'b0000101000010100010 : color = 12'he73;
15'b0000101000010100011 : color = 12'he73;
15'b0000101000010100100 : color = 12'he73;
15'b0000101000010100101 : color = 12'he73;
15'b0000101000010100110 : color = 12'he73;
15'b0000101000010100111 : color = 12'he73;
15'b0000101000010101000 : color = 12'he73;
15'b0000101000010101001 : color = 12'he51;
15'b0000101000010101010 : color = 12'hf00;
15'b0000101000010101011 : color = 12'hf11;
15'b0000101000010101100 : color = 12'hf73;
15'b0000101000010101101 : color = 12'he73;
15'b0000101000010101110 : color = 12'he73;
15'b0000101000010101111 : color = 12'he73;
15'b0000101000010110000 : color = 12'he73;
15'b0000101000010110001 : color = 12'he73;
15'b0000101000010110010 : color = 12'he73;
15'b0000101000010110011 : color = 12'he61;
15'b0000101000010110100 : color = 12'hf31;
15'b0000101000010110101 : color = 12'hf52;
15'b0000101000010110110 : color = 12'hf73;
15'b0000101000010110111 : color = 12'he73;
15'b0000101000010111000 : color = 12'hf51;
15'b0000101000010111001 : color = 12'hf31;
15'b0000101000010111010 : color = 12'hf63;
15'b0000101000010111011 : color = 12'he73;
15'b0000101000010111100 : color = 12'he73;
15'b0000101000010111101 : color = 12'he73;
15'b0000101000010111110 : color = 12'he73;
15'b0000101000010111111 : color = 12'he73;
15'b0000101000011000000 : color = 12'he73;
15'b0000101000011000001 : color = 12'he73;
15'b0000101000011000010 : color = 12'he73;
15'b0000101000011000011 : color = 12'he73;
15'b0000101000011000100 : color = 12'he73;
15'b0000101000011000101 : color = 12'he73;
15'b0000101000011000110 : color = 12'he73;
15'b0000101000011000111 : color = 12'he73;
15'b0000101000011001000 : color = 12'he73;
15'b0000101000011001001 : color = 12'he73;
15'b0000101000011001010 : color = 12'he73;
15'b0000101000011001011 : color = 12'he73;
15'b0000101000011001100 : color = 12'he73;
15'b0000101000011001101 : color = 12'he73;
15'b0000101000011001110 : color = 12'he73;
15'b0000101000011001111 : color = 12'he73;
15'b0000101000011010000 : color = 12'he73;
15'b0000101000011010001 : color = 12'he73;
15'b0000101000011010010 : color = 12'he73;
15'b0000101000011010011 : color = 12'he73;
15'b0000101000011010100 : color = 12'he73;
15'b0000101000011010101 : color = 12'he73;
15'b0000101000011010110 : color = 12'he73;
15'b0000101000011010111 : color = 12'hf30;
15'b0000101000011011000 : color = 12'hf01;
15'b0000101000011011001 : color = 12'hf73;
15'b0000101000011011010 : color = 12'he73;
15'b0000101000011011011 : color = 12'he73;
15'b0000101000011011100 : color = 12'he62;
15'b0000101000011011101 : color = 12'hf31;
15'b0000101000011011110 : color = 12'hf31;
15'b0000101000011011111 : color = 12'hf31;
15'b0000101000011100000 : color = 12'hf31;
15'b0000101000011100001 : color = 12'hf31;
15'b0000101000011100010 : color = 12'hf31;
15'b0000101000011100011 : color = 12'hf31;
15'b0000101000011100100 : color = 12'hf31;
15'b0000101000011100101 : color = 12'hf31;
15'b0000101000011100110 : color = 12'hf31;
15'b0000101000011100111 : color = 12'hf31;
15'b0000101000011101000 : color = 12'hf30;
15'b0000101000011101001 : color = 12'hf00;
15'b0000101000011101010 : color = 12'hf00;
15'b0000101000011101011 : color = 12'hf11;
15'b0000101000011101100 : color = 12'hf73;
15'b0000101000011101101 : color = 12'he73;
15'b0000101000011101110 : color = 12'he73;
15'b0000101000011101111 : color = 12'he73;
15'b0000101000011110000 : color = 12'he73;
15'b0000101000011110001 : color = 12'he73;
15'b0000101000011110010 : color = 12'he73;
15'b0000101000011110011 : color = 12'he73;
15'b0000101000011110100 : color = 12'he73;
15'b0000101000011110101 : color = 12'he73;
15'b0000101000011110110 : color = 12'he73;
15'b0000101000011110111 : color = 12'he73;
15'b0000101000011111000 : color = 12'he73;
15'b0000101000011111001 : color = 12'he73;
15'b0000101000011111010 : color = 12'he73;
15'b0000101000011111011 : color = 12'he73;
15'b0000101000011111100 : color = 12'he73;
15'b0000101000011111101 : color = 12'he73;
15'b0000101000011111110 : color = 12'he73;
15'b0000101000011111111 : color = 12'he73;
15'b0000101000100000000 : color = 12'he73;
15'b0000101000100000001 : color = 12'hf30;
15'b0000101000100000010 : color = 12'hf11;
15'b0000101000100000011 : color = 12'hf73;
15'b0000101000100000100 : color = 12'he73;
15'b0000101000100000101 : color = 12'hf31;
15'b0000101000100000110 : color = 12'hf63;
15'b0000101000100000111 : color = 12'he73;
15'b0000101000100001000 : color = 12'he73;
15'b0000101000100001001 : color = 12'he73;
15'b0000101000100001010 : color = 12'he73;
15'b0000101000100001011 : color = 12'he73;
15'b0000101000100001100 : color = 12'hf40;
15'b0000101000100001101 : color = 12'hf32;
15'b0000101000100001110 : color = 12'hf73;
15'b0000101000100001111 : color = 12'he73;
15'b0000101000100010000 : color = 12'he51;
15'b0000101000100010001 : color = 12'hf32;
15'b0000101000100010010 : color = 12'hf73;
15'b0000101000100010011 : color = 12'he73;
15'b0000101000100010100 : color = 12'he73;
15'b0000101000100010101 : color = 12'he73;
15'b0000101000100010110 : color = 12'he73;
15'b0000101000100010111 : color = 12'he73;
15'b0000101000100011000 : color = 12'he73;
15'b0000101000100011001 : color = 12'he73;
15'b0000101000100011010 : color = 12'he73;
15'b0000101000100011011 : color = 12'he73;
15'b0000101000100011100 : color = 12'he73;
15'b0000101000100011101 : color = 12'he73;
15'b0000101000100011110 : color = 12'he73;
15'b0000101000100011111 : color = 12'he73;
15'b0000101000100100000 : color = 12'he73;
15'b0000101000100100001 : color = 12'he73;
15'b0000101000100100010 : color = 12'he73;
15'b0000101000100100011 : color = 12'he73;
15'b0000101000100100100 : color = 12'he73;
15'b0000101000100100101 : color = 12'he73;
15'b0000101000100100110 : color = 12'he73;
15'b0000101000100100111 : color = 12'he73;
15'b0000101000100101000 : color = 12'he73;
15'b0000101000100101001 : color = 12'he73;
15'b0000101000100101010 : color = 12'he72;
15'b0000101000100101011 : color = 12'hf31;
15'b0000101000100101100 : color = 12'hf31;
15'b0000101000100101101 : color = 12'hf31;
15'b0000101000100101110 : color = 12'hf31;
15'b0000101000100101111 : color = 12'hf31;
15'b0000101000100110000 : color = 12'hf31;
15'b0000101000100110001 : color = 12'hf30;
15'b0000101000100110010 : color = 12'hf00;
15'b0000101000100110011 : color = 12'hf00;
15'b0000101000100110100 : color = 12'hf42;
15'b0000101000100110101 : color = 12'he61;
15'b0000101000100110110 : color = 12'hf00;
15'b0000101000100110111 : color = 12'hf63;
15'b0000101000100111000 : color = 12'he73;
15'b0000101000100111001 : color = 12'he73;
15'b0000101000100111010 : color = 12'he73;
15'b0000101000100111011 : color = 12'hf30;
15'b0000101000100111100 : color = 12'hf32;
15'b0000101000100111101 : color = 12'he73;
15'b0000101000100111110 : color = 12'he73;
15'b0000101000100111111 : color = 12'he73;
15'b0000101000101000000 : color = 12'he61;
15'b0000101000101000001 : color = 12'hf00;
15'b0000101000101000010 : color = 12'hf63;
15'b0000101000101000011 : color = 12'he73;
15'b0000101000101000100 : color = 12'he73;
15'b0000101000101000101 : color = 12'he73;
15'b0000101000101000110 : color = 12'he73;
15'b0000101000101000111 : color = 12'he73;
15'b0000101000101001000 : color = 12'he73;
15'b0000101000101001001 : color = 12'he73;
15'b0000101000101001010 : color = 12'he73;
15'b0000101000101001011 : color = 12'he73;
15'b0000101000101001100 : color = 12'he73;
15'b0000101000101001101 : color = 12'he73;
15'b0000101000101001110 : color = 12'he73;
15'b0000101000101001111 : color = 12'he73;
15'b0000101000101010000 : color = 12'he73;
15'b0000101000101010001 : color = 12'he73;
15'b0000101000101010010 : color = 12'he73;
15'b0000101000101010011 : color = 12'he73;
15'b0000101000101010100 : color = 12'he73;
15'b0000101000101010101 : color = 12'he73;
15'b0000101000101010110 : color = 12'he73;
15'b0000101000101010111 : color = 12'he73;
15'b0000101000101011000 : color = 12'he73;
15'b0000101000101011001 : color = 12'he73;
15'b0000101000101011010 : color = 12'he73;
15'b0000101000101011011 : color = 12'he73;
15'b0000101000101011100 : color = 12'he73;
15'b0000101000101011101 : color = 12'he73;
15'b0000101000101011110 : color = 12'he73;
15'b0000101000101011111 : color = 12'he73;
15'b0000101000101100000 : color = 12'he73;
15'b0000101000101100001 : color = 12'he72;
15'b0000101000101100010 : color = 12'hf00;
15'b0000101000101100011 : color = 12'hf00;
15'b0000101000101100100 : color = 12'hf31;
15'b0000101000101100101 : color = 12'hf63;
15'b0000101000101100110 : color = 12'he73;
15'b0000101000101100111 : color = 12'he73;
15'b0000101000101101000 : color = 12'he73;
15'b0000101000101101001 : color = 12'he73;
15'b0000101000101101010 : color = 12'he73;
15'b0000101000101101011 : color = 12'he73;
15'b0000101000101101100 : color = 12'he73;
15'b0000101000101101101 : color = 12'he73;
15'b0000101000101101110 : color = 12'he73;
15'b0000101000101101111 : color = 12'he73;
15'b0000101000101110000 : color = 12'he73;
15'b0000101000101110001 : color = 12'he73;
15'b0000101000101110010 : color = 12'he73;
15'b0000101000101110011 : color = 12'he73;
15'b0000101000101110100 : color = 12'he73;
15'b0000101000101110101 : color = 12'he73;
15'b0000101000101110110 : color = 12'he73;
15'b0000101000101110111 : color = 12'he73;
15'b0000101000101111000 : color = 12'he73;
15'b0000101000101111001 : color = 12'he73;
15'b0000101000101111010 : color = 12'he73;
15'b0000101000101111011 : color = 12'he73;
15'b0000101000101111100 : color = 12'he73;
15'b0000101000101111101 : color = 12'he73;
15'b0000101000101111110 : color = 12'he73;
15'b0000101000101111111 : color = 12'he73;
15'b0000101000110000000 : color = 12'he73;
15'b0000101000110000001 : color = 12'he73;
15'b0000101000110000010 : color = 12'he73;
15'b0000101000110000011 : color = 12'he73;
15'b0000101000110000100 : color = 12'he73;
15'b0000101000110000101 : color = 12'he73;
15'b0000101000110000110 : color = 12'he51;
15'b0000101000110000111 : color = 12'hf00;
15'b0000101000110001000 : color = 12'hf63;
15'b0000101000110001001 : color = 12'he73;
15'b0000101000110001010 : color = 12'he73;
15'b0000101000110001011 : color = 12'he73;
15'b0000101000110001100 : color = 12'he62;
15'b0000101000110001101 : color = 12'hf31;
15'b0000101000110001110 : color = 12'hf31;
15'b0000101000110001111 : color = 12'hf31;
15'b0000101000110010000 : color = 12'hf31;
15'b0000101000110010001 : color = 12'hf31;
15'b0000101000110010010 : color = 12'hf31;
15'b0000101000110010011 : color = 12'hf10;
15'b0000101000110010100 : color = 12'hf11;
15'b0000101000110010101 : color = 12'hf31;
15'b0000101000110010110 : color = 12'hf31;
15'b0000101000110010111 : color = 12'hf31;
15'b0000101000110011000 : color = 12'hf30;
15'b0000101000110011001 : color = 12'hf00;
15'b0000101000110011010 : color = 12'hf00;
15'b0000101000110011011 : color = 12'hf11;
15'b0000101000110011100 : color = 12'hf73;
15'b0000101000110011101 : color = 12'he73;
15'b0000101000110011110 : color = 12'he73;
15'b0000101000110011111 : color = 12'he73;
15'b0000101000110100000 : color = 12'he73;
15'b0000101000110100001 : color = 12'he73;
15'b0000101000110100010 : color = 12'he73;
15'b0000101000110100011 : color = 12'he73;
15'b0000101000110100100 : color = 12'he73;
15'b0000101000110100101 : color = 12'he73;
15'b0000101000110100110 : color = 12'he73;
15'b0000101000110100111 : color = 12'he73;
15'b0000101000110101000 : color = 12'he73;
15'b0000101000110101001 : color = 12'he73;
15'b0000101000110101010 : color = 12'he73;
15'b0000101000110101011 : color = 12'he73;
15'b0000101000110101100 : color = 12'he73;
15'b0000100111111101011 : color = 12'he73;
15'b0000100111111101100 : color = 12'he73;
15'b0000100111111101101 : color = 12'he73;
15'b0000100111111101110 : color = 12'he73;
15'b0000100111111101111 : color = 12'he73;
15'b0000100111111110000 : color = 12'he73;
15'b0000100111111110001 : color = 12'he73;
15'b0000100111111110010 : color = 12'he73;
15'b0000100111111110011 : color = 12'he73;
15'b0000100111111110100 : color = 12'he73;
15'b0000100111111110101 : color = 12'he73;
15'b0000100111111110110 : color = 12'he73;
15'b0000100111111110111 : color = 12'he73;
15'b0000100111111111000 : color = 12'he73;
15'b0000100111111111001 : color = 12'he73;
15'b0000100111111111010 : color = 12'he73;
15'b0000100111111111011 : color = 12'he72;
15'b0000100111111111100 : color = 12'hf00;
15'b0000100111111111101 : color = 12'hf31;
15'b0000100111111111110 : color = 12'hf73;
15'b0000100111111111111 : color = 12'he73;
15'b0000101000000000000 : color = 12'he73;
15'b0000101000000000001 : color = 12'he51;
15'b0000101000000000010 : color = 12'hf00;
15'b0000101000000000011 : color = 12'hf53;
15'b0000101000000000100 : color = 12'he73;
15'b0000101000000000101 : color = 12'he73;
15'b0000101000000000110 : color = 12'he73;
15'b0000101000000000111 : color = 12'he73;
15'b0000101000000001000 : color = 12'he73;
15'b0000101000000001001 : color = 12'he73;
15'b0000101000000001010 : color = 12'he73;
15'b0000101000000001011 : color = 12'he73;
15'b0000101000000001100 : color = 12'he73;
15'b0000101000000001101 : color = 12'he73;
15'b0000101000000001110 : color = 12'he73;
15'b0000101000000001111 : color = 12'he73;
15'b0000101000000010000 : color = 12'he73;
15'b0000101000000010001 : color = 12'he73;
15'b0000101000000010010 : color = 12'he73;
15'b0000101000000010011 : color = 12'he73;
15'b0000101000000010100 : color = 12'he73;
15'b0000101000000010101 : color = 12'he73;
15'b0000101000000010110 : color = 12'he73;
15'b0000101000000010111 : color = 12'he73;
15'b0000101000000011000 : color = 12'he73;
15'b0000101000000011001 : color = 12'he73;
15'b0000101000000011010 : color = 12'he73;
15'b0000101000000011011 : color = 12'he73;
15'b0000101000000011100 : color = 12'he73;
15'b0000101000000011101 : color = 12'he73;
15'b0000101000000011110 : color = 12'he73;
15'b0000101000000011111 : color = 12'he73;
15'b0000101000000100000 : color = 12'he73;
15'b0000101000000100001 : color = 12'he73;
15'b0000101000000100010 : color = 12'he73;
15'b0000101000000100011 : color = 12'he51;
15'b0000101000000100100 : color = 12'hf00;
15'b0000101000000100101 : color = 12'hf42;
15'b0000101000000100110 : color = 12'he73;
15'b0000101000000100111 : color = 12'he73;
15'b0000101000000101000 : color = 12'he61;
15'b0000101000000101001 : color = 12'hf00;
15'b0000101000000101010 : color = 12'hf53;
15'b0000101000000101011 : color = 12'he73;
15'b0000101000000101100 : color = 12'he73;
15'b0000101000000101101 : color = 12'he73;
15'b0000101000000101110 : color = 12'he73;
15'b0000101000000101111 : color = 12'he72;
15'b0000101000000110000 : color = 12'hf00;
15'b0000101000000110001 : color = 12'hf11;
15'b0000101000000110010 : color = 12'hf31;
15'b0000101000000110011 : color = 12'hf31;
15'b0000101000000110100 : color = 12'hf31;
15'b0000101000000110101 : color = 12'hf31;
15'b0000101000000110110 : color = 12'hf00;
15'b0000101000000110111 : color = 12'hf00;
15'b0000101000000111000 : color = 12'hf53;
15'b0000101000000111001 : color = 12'he73;
15'b0000101000000111010 : color = 12'he73;
15'b0000101000000111011 : color = 12'he73;
15'b0000101000000111100 : color = 12'he73;
15'b0000101000000111101 : color = 12'he73;
15'b0000101000000111110 : color = 12'he73;
15'b0000101000000111111 : color = 12'he73;
15'b0000101000001000000 : color = 12'he73;
15'b0000101000001000001 : color = 12'he73;
15'b0000101000001000010 : color = 12'he73;
15'b0000101000001000011 : color = 12'he73;
15'b0000101000001000100 : color = 12'he73;
15'b0000101000001000101 : color = 12'he73;
15'b0000101000001000110 : color = 12'he73;
15'b0000101000001000111 : color = 12'he73;
15'b0000101000001001000 : color = 12'he73;
15'b0000101000001001001 : color = 12'he73;
15'b0000101000001001010 : color = 12'he73;
15'b0000101000001001011 : color = 12'he73;
15'b0000101000001001100 : color = 12'he73;
15'b0000101000001001101 : color = 12'he62;
15'b0000101000001001110 : color = 12'hf31;
15'b0000101000001001111 : color = 12'hf31;
15'b0000101000001010000 : color = 12'hf31;
15'b0000101000001010001 : color = 12'hf31;
15'b0000101000001010010 : color = 12'hf31;
15'b0000101000001010011 : color = 12'hf31;
15'b0000101000001010100 : color = 12'hf31;
15'b0000101000001010101 : color = 12'hf31;
15'b0000101000001010110 : color = 12'hf31;
15'b0000101000001010111 : color = 12'hf10;
15'b0000101000001011000 : color = 12'hf00;
15'b0000101000001011001 : color = 12'hf11;
15'b0000101000001011010 : color = 12'hf31;
15'b0000101000001011011 : color = 12'hf31;
15'b0000101000001011100 : color = 12'hf31;
15'b0000101000001011101 : color = 12'hf31;
15'b0000101000001011110 : color = 12'hf31;
15'b0000101000001011111 : color = 12'hf31;
15'b0000101000001100000 : color = 12'hf10;
15'b0000101000001100001 : color = 12'hf00;
15'b0000101000001100010 : color = 12'hf00;
15'b0000101000001100011 : color = 12'hf42;
15'b0000101000001100100 : color = 12'he73;
15'b0000101000001100101 : color = 12'he73;
15'b0000101000001100110 : color = 12'he73;
15'b0000101000001100111 : color = 12'he73;
15'b0000101000001101000 : color = 12'he73;
15'b0000101000001101001 : color = 12'he73;
15'b0000101000001101010 : color = 12'he73;
15'b0000101000001101011 : color = 12'he73;
15'b0000101000001101100 : color = 12'he73;
15'b0000101000001101101 : color = 12'he73;
15'b0000101000001101110 : color = 12'he73;
15'b0000101000001101111 : color = 12'he73;
15'b0000101000001110000 : color = 12'he73;
15'b0000101000001110001 : color = 12'he73;
15'b0000101000001110010 : color = 12'he73;
15'b0000101000001110011 : color = 12'he73;
15'b0000101000001110100 : color = 12'he73;
15'b0000101000001110101 : color = 12'he73;
15'b0000101000001110110 : color = 12'he73;
15'b0000101000001110111 : color = 12'he73;
15'b0000101000001111000 : color = 12'he73;
15'b0000101000001111001 : color = 12'he73;
15'b0000101000001111010 : color = 12'he73;
15'b0000101000001111011 : color = 12'he73;
15'b0000101000001111100 : color = 12'he73;
15'b0000101000001111101 : color = 12'he73;
15'b0000101000001111110 : color = 12'hf30;
15'b0000101000001111111 : color = 12'hf00;
15'b0000101000010000000 : color = 12'hf31;
15'b0000101000010000001 : color = 12'hf63;
15'b0000101000010000010 : color = 12'he73;
15'b0000101000010000011 : color = 12'he73;
15'b0000101000010000100 : color = 12'he73;
15'b0000101000010000101 : color = 12'he73;
15'b0000101000010000110 : color = 12'he73;
15'b0000101000010000111 : color = 12'he73;
15'b0000101000010001000 : color = 12'he72;
15'b0000101000010001001 : color = 12'hf00;
15'b0000101000010001010 : color = 12'hf52;
15'b0000101000010001011 : color = 12'hf73;
15'b0000101000010001100 : color = 12'he73;
15'b0000101000010001101 : color = 12'he73;
15'b0000101000010001110 : color = 12'hf40;
15'b0000101000010001111 : color = 12'hf01;
15'b0000101000010010000 : color = 12'hf73;
15'b0000101000010010001 : color = 12'he73;
15'b0000101000010010010 : color = 12'he73;
15'b0000101000010010011 : color = 12'he73;
15'b0000101000010010100 : color = 12'he73;
15'b0000101000010010101 : color = 12'he73;
15'b0000101000010010110 : color = 12'he73;
15'b0000101000010010111 : color = 12'he73;
15'b0000101000010011000 : color = 12'he73;
15'b0000101000010011001 : color = 12'he73;
15'b0000101000010011010 : color = 12'he73;
15'b0000101000010011011 : color = 12'he73;
15'b0000101000010011100 : color = 12'he73;
15'b0000101000010011101 : color = 12'he73;
15'b0000101000010011110 : color = 12'he73;
15'b0000101000010011111 : color = 12'he73;
15'b0000101000010100000 : color = 12'he73;
15'b0000101000010100001 : color = 12'he73;
15'b0000101000010100010 : color = 12'he73;
15'b0000101000010100011 : color = 12'he72;
15'b0000101000010100100 : color = 12'hf41;
15'b0000101000010100101 : color = 12'hf31;
15'b0000101000010100110 : color = 12'hf31;
15'b0000101000010100111 : color = 12'hf31;
15'b0000101000010101000 : color = 12'hf31;
15'b0000101000010101001 : color = 12'hf31;
15'b0000101000010101010 : color = 12'hf31;
15'b0000101000010101011 : color = 12'hf31;
15'b0000101000010101100 : color = 12'hf31;
15'b0000101000010101101 : color = 12'hf31;
15'b0000101000010101110 : color = 12'hf31;
15'b0000101000010101111 : color = 12'hf31;
15'b0000101000010110000 : color = 12'hf31;
15'b0000101000010110001 : color = 12'hf31;
15'b0000101000010110010 : color = 12'hf31;
15'b0000101000010110011 : color = 12'hf31;
15'b0000101000010110100 : color = 12'hf31;
15'b0000101000010110101 : color = 12'hf31;
15'b0000101000010110110 : color = 12'hf31;
15'b0000101000010110111 : color = 12'hf31;
15'b0000101000010111000 : color = 12'hf31;
15'b0000101000010111001 : color = 12'hf00;
15'b0000101000010111010 : color = 12'hf00;
15'b0000101000010111011 : color = 12'hf00;
15'b0000101000010111100 : color = 12'hf11;
15'b0000101000010111101 : color = 12'hf73;
15'b0000101000010111110 : color = 12'he73;
15'b0000101000010111111 : color = 12'he73;
15'b0000101000011000000 : color = 12'he73;
15'b0000101000011000001 : color = 12'he73;
15'b0000101000011000010 : color = 12'he73;
15'b0000101000011000011 : color = 12'he73;
15'b0000101000011000100 : color = 12'he73;
15'b0000101000011000101 : color = 12'he73;
15'b0000101000011000110 : color = 12'he73;
15'b0000101000011000111 : color = 12'he73;
15'b0000101000011001000 : color = 12'he73;
15'b0000101000011001001 : color = 12'he73;
15'b0000101000011001010 : color = 12'he73;
15'b0000101000011001011 : color = 12'he73;
15'b0000101000011001100 : color = 12'he73;
15'b0000101000011001101 : color = 12'he73;
15'b0000101000011001110 : color = 12'he73;
15'b0000101000011001111 : color = 12'he73;
15'b0000101000011010000 : color = 12'he73;
15'b0000101000011010001 : color = 12'he73;
15'b0000101000011010010 : color = 12'he72;
15'b0000101000011010011 : color = 12'hf10;
15'b0000101000011010100 : color = 12'hf01;
15'b0000101000011010101 : color = 12'hf73;
15'b0000101000011010110 : color = 12'he73;
15'b0000101000011010111 : color = 12'he73;
15'b0000101000011011000 : color = 12'he73;
15'b0000101000011011001 : color = 12'he73;
15'b0000101000011011010 : color = 12'he73;
15'b0000101000011011011 : color = 12'he73;
15'b0000101000011011100 : color = 12'he73;
15'b0000101000011011101 : color = 12'he62;
15'b0000101000011011110 : color = 12'hf10;
15'b0000101000011011111 : color = 12'hf00;
15'b0000101000011100000 : color = 12'hf31;
15'b0000101000011100001 : color = 12'hf63;
15'b0000101000011100010 : color = 12'he73;
15'b0000101000011100011 : color = 12'he73;
15'b0000101000011100100 : color = 12'he73;
15'b0000101000011100101 : color = 12'he73;
15'b0000101000011100110 : color = 12'he73;
15'b0000101000011100111 : color = 12'he73;
15'b0000101000011101000 : color = 12'he73;
15'b0000101000011101001 : color = 12'he73;
15'b0000101000011101010 : color = 12'he73;
15'b0000101000011101011 : color = 12'he73;
15'b0000101000011101100 : color = 12'he73;
15'b0000101000011101101 : color = 12'he73;
15'b0000101000011101110 : color = 12'he73;
15'b0000101000011101111 : color = 12'he73;
15'b0000101000011110000 : color = 12'he73;
15'b0000101000011110001 : color = 12'he73;
15'b0000101000011110010 : color = 12'he73;
15'b0000101000011110011 : color = 12'he73;
15'b0000101000011110100 : color = 12'he73;
15'b0000101000011110101 : color = 12'he73;
15'b0000101000011110110 : color = 12'he73;
15'b0000101000011110111 : color = 12'he73;
15'b0000101000011111000 : color = 12'he73;
15'b0000101000011111001 : color = 12'he73;
15'b0000101000011111010 : color = 12'he73;
15'b0000101000011111011 : color = 12'he73;
15'b0000101000011111100 : color = 12'he73;
15'b0000101000011111101 : color = 12'he73;
15'b0000101000011111110 : color = 12'he73;
15'b0000101000011111111 : color = 12'he73;
15'b0000101000100000000 : color = 12'hf40;
15'b0000101000100000001 : color = 12'hf01;
15'b0000101000100000010 : color = 12'hf73;
15'b0000101000100000011 : color = 12'he73;
15'b0000101000100000100 : color = 12'he73;
15'b0000101000100000101 : color = 12'he73;
15'b0000101000100000110 : color = 12'he62;
15'b0000101000100000111 : color = 12'hf63;
15'b0000101000100001000 : color = 12'he73;
15'b0000101000100001001 : color = 12'he73;
15'b0000101000100001010 : color = 12'he73;
15'b0000101000100001011 : color = 12'he73;
15'b0000101000100001100 : color = 12'he51;
15'b0000101000100001101 : color = 12'hf00;
15'b0000101000100001110 : color = 12'hf53;
15'b0000101000100001111 : color = 12'he73;
15'b0000101000100010000 : color = 12'he73;
15'b0000101000100010001 : color = 12'he73;
15'b0000101000100010010 : color = 12'he73;
15'b0000101000100010011 : color = 12'he73;
15'b0000101000100010100 : color = 12'he73;
15'b0000101000100010101 : color = 12'he73;
15'b0000101000100010110 : color = 12'he73;
15'b0000101000100010111 : color = 12'he73;
15'b0000101000100011000 : color = 12'he73;
15'b0000101000100011001 : color = 12'he73;
15'b0000101000100011010 : color = 12'he73;
15'b0000101000100011011 : color = 12'he73;
15'b0000101000100011100 : color = 12'he73;
15'b0000101000100011101 : color = 12'he73;
15'b0000101000100011110 : color = 12'he73;
15'b0000101000100011111 : color = 12'he73;
15'b0000101000100100000 : color = 12'he73;
15'b0000101000100100001 : color = 12'he73;
15'b0000101000100100010 : color = 12'he73;
15'b0000101000100100011 : color = 12'he73;
15'b0000101000100100100 : color = 12'he73;
15'b0000101000100100101 : color = 12'he73;
15'b0000101000100100110 : color = 12'he73;
15'b0000101000100100111 : color = 12'he73;
15'b0000101000100101000 : color = 12'he73;
15'b0000101000100101001 : color = 12'he51;
15'b0000101000100101010 : color = 12'hf11;
15'b0000101000100101011 : color = 12'hf73;
15'b0000101000100101100 : color = 12'he73;
15'b0000101000100101101 : color = 12'he73;
15'b0000101000100101110 : color = 12'he51;
15'b0000101000100101111 : color = 12'hf00;
15'b0000101000100110000 : color = 12'hf63;
15'b0000101000100110001 : color = 12'he73;
15'b0000101000100110010 : color = 12'he73;
15'b0000101000100110011 : color = 12'he73;
15'b0000101000100110100 : color = 12'he51;
15'b0000101000100110101 : color = 12'hf52;
15'b0000101000100110110 : color = 12'he73;
15'b0000101000100110111 : color = 12'he73;
15'b0000101000100111000 : color = 12'he73;
15'b0000101000100111001 : color = 12'he73;
15'b0000101000100111010 : color = 12'hf30;
15'b0000101000100111011 : color = 12'hf11;
15'b0000101000100111100 : color = 12'hf73;
15'b0000101000100111101 : color = 12'he73;
15'b0000101000100111110 : color = 12'he73;
15'b0000101000100111111 : color = 12'he73;
15'b0000101000101000000 : color = 12'he73;
15'b0000101000101000001 : color = 12'he73;
15'b0000101000101000010 : color = 12'he73;
15'b0000101000101000011 : color = 12'he73;
15'b0000101000101000100 : color = 12'he73;
15'b0000101000101000101 : color = 12'he73;
15'b0000101000101000110 : color = 12'he73;
15'b0000101000101000111 : color = 12'he73;
15'b0000101000101001000 : color = 12'he73;
15'b0000101000101001001 : color = 12'he73;
15'b0000101000101001010 : color = 12'he73;
15'b0000101000101001011 : color = 12'he73;
15'b0000101000101001100 : color = 12'he73;
15'b0000101000101001101 : color = 12'he73;
15'b0000101000101001110 : color = 12'he73;
15'b0000101000101001111 : color = 12'he73;
15'b0000101000101010000 : color = 12'he73;
15'b0000101000101010001 : color = 12'he73;
15'b0000101000101010010 : color = 12'he73;
15'b0000101000101010011 : color = 12'he73;
15'b0000101000101010100 : color = 12'he62;
15'b0000101000101010101 : color = 12'hf63;
15'b0000101000101010110 : color = 12'he73;
15'b0000101000101010111 : color = 12'he72;
15'b0000101000101011000 : color = 12'hf10;
15'b0000101000101011001 : color = 12'hf32;
15'b0000101000101011010 : color = 12'he73;
15'b0000101000101011011 : color = 12'he73;
15'b0000101000101011100 : color = 12'he73;
15'b0000101000101011101 : color = 12'he73;
15'b0000101000101011110 : color = 12'he61;
15'b0000101000101011111 : color = 12'hf00;
15'b0000101000101100000 : color = 12'hf63;
15'b0000101000101100001 : color = 12'he73;
15'b0000101000101100010 : color = 12'he73;
15'b0000101000101100011 : color = 12'he73;
15'b0000101000101100100 : color = 12'hf30;
15'b0000101000101100101 : color = 12'hf32;
15'b0000101000101100110 : color = 12'he73;
15'b0000101000101100111 : color = 12'he73;
15'b0000101000101101000 : color = 12'he73;
15'b0000101000101101001 : color = 12'he61;
15'b0000101000101101010 : color = 12'hf00;
15'b0000101000101101011 : color = 12'hf63;
15'b0000101000101101100 : color = 12'he73;
15'b0000101000101101101 : color = 12'he73;
15'b0000101000101101110 : color = 12'he73;
15'b0000101000101101111 : color = 12'he73;
15'b0000101000101110000 : color = 12'he73;
15'b0000101000101110001 : color = 12'he73;
15'b0000101000101110010 : color = 12'he73;
15'b0000101000101110011 : color = 12'he73;
15'b0000101000101110100 : color = 12'he73;
15'b0000101000101110101 : color = 12'he73;
15'b0000101000101110110 : color = 12'he73;
15'b0000101000101110111 : color = 12'he73;
15'b0000101000101111000 : color = 12'he73;
15'b0000101000101111001 : color = 12'he73;
15'b0000101000101111010 : color = 12'he73;
15'b0000101000101111011 : color = 12'he73;
15'b0000101000101111100 : color = 12'he73;
15'b0000101000101111101 : color = 12'he73;
15'b0000101000101111110 : color = 12'he73;
15'b0000101000101111111 : color = 12'he73;
15'b0000101000110000000 : color = 12'he73;
15'b0000101000110000001 : color = 12'he73;
15'b0000101000110000010 : color = 12'he73;
15'b0000101000110000011 : color = 12'he73;
15'b0000101000110000100 : color = 12'he73;
15'b0000101000110000101 : color = 12'he73;
15'b0000101000110000110 : color = 12'he73;
15'b0000101000110000111 : color = 12'he73;
15'b0000101000110001000 : color = 12'he73;
15'b0000101000110001001 : color = 12'he72;
15'b0000101000110001010 : color = 12'hf10;
15'b0000101000110001011 : color = 12'hf11;
15'b0000101000110001100 : color = 12'hf63;
15'b0000101000110001101 : color = 12'he73;
15'b0000101000110001110 : color = 12'he73;
15'b0000101000110001111 : color = 12'he73;
15'b0000101000110010000 : color = 12'he73;
15'b0000101000110010001 : color = 12'he73;
15'b0000101000110010010 : color = 12'he73;
15'b0000101000110010011 : color = 12'he73;
15'b0000101000110010100 : color = 12'he73;
15'b0000101000110010101 : color = 12'he73;
15'b0000101000110010110 : color = 12'he73;
15'b0000101000110010111 : color = 12'he73;
15'b0000101000110011000 : color = 12'he73;
15'b0000101000110011001 : color = 12'he73;
15'b0000101000110011010 : color = 12'he73;
15'b0000101000110011011 : color = 12'he73;
15'b0000101000110011100 : color = 12'he73;
15'b0000101000110011101 : color = 12'he73;
15'b0000101000110011110 : color = 12'he73;
15'b0000101000110011111 : color = 12'he73;
15'b0000101000110100000 : color = 12'he73;
15'b0000101000110100001 : color = 12'he73;
15'b0000101000110100010 : color = 12'he73;
15'b0000101000110100011 : color = 12'he73;
15'b0000101000110100100 : color = 12'he73;
15'b0000101000110100101 : color = 12'he73;
15'b0000101000110100110 : color = 12'he73;
15'b0000101000110100111 : color = 12'he73;
15'b0000101000110101000 : color = 12'he73;
15'b0000101000110101001 : color = 12'he73;
15'b0000101000110101010 : color = 12'he73;
15'b0000101000110101011 : color = 12'he73;
15'b0000101000110101100 : color = 12'he73;
15'b0000101000110101101 : color = 12'he73;
15'b0000101000110101110 : color = 12'he72;
15'b0000101000110101111 : color = 12'hf10;
15'b0000101000110110000 : color = 12'hf42;
15'b0000101000110110001 : color = 12'he73;
15'b0000101000110110010 : color = 12'he73;
15'b0000101000110110011 : color = 12'he73;
15'b0000101000110110100 : color = 12'hf62;
15'b0000101000110110101 : color = 12'he73;
15'b0000101000110110110 : color = 12'hf62;
15'b0000101000110110111 : color = 12'hf73;
15'b0000101000110111000 : color = 12'he73;
15'b0000101000110111001 : color = 12'he73;
15'b0000101000110111010 : color = 12'he73;
15'b0000101000110111011 : color = 12'hf40;
15'b0000101000110111100 : color = 12'hf11;
15'b0000101000110111101 : color = 12'hf73;
15'b0000101000110111110 : color = 12'he73;
15'b0000101000110111111 : color = 12'he73;
15'b0000101000111000000 : color = 12'he73;
15'b0000101000111000001 : color = 12'he73;
15'b0000101000111000010 : color = 12'he73;
15'b0000101000111000011 : color = 12'he73;
15'b0000101000111000100 : color = 12'he73;
15'b0000101000111000101 : color = 12'he73;
15'b0000101000111000110 : color = 12'he73;
15'b0000101000111000111 : color = 12'he73;
15'b0000101000111001000 : color = 12'he73;
15'b0000101000111001001 : color = 12'he73;
15'b0000101000111001010 : color = 12'he73;
15'b0000101000111001011 : color = 12'he73;
15'b0000101000111001100 : color = 12'he73;
15'b0000101000111001101 : color = 12'he73;
15'b0000101000111001110 : color = 12'he73;
15'b0000101000111001111 : color = 12'he73;
15'b0000101000111010000 : color = 12'he73;
15'b0000101000111010001 : color = 12'he73;
15'b0000101000111010010 : color = 12'he73;
15'b0000101000111010011 : color = 12'he73;
15'b0000101000111010100 : color = 12'he73;
15'b0000101000111010101 : color = 12'he73;
15'b0000101000000010100 : color = 12'he73;
15'b0000101000000010101 : color = 12'he73;
15'b0000101000000010110 : color = 12'he73;
15'b0000101000000010111 : color = 12'he73;
15'b0000101000000011000 : color = 12'he73;
15'b0000101000000011001 : color = 12'he73;
15'b0000101000000011010 : color = 12'he73;
15'b0000101000000011011 : color = 12'he73;
15'b0000101000000011100 : color = 12'he73;
15'b0000101000000011101 : color = 12'he73;
15'b0000101000000011110 : color = 12'he73;
15'b0000101000000011111 : color = 12'he73;
15'b0000101000000100000 : color = 12'he73;
15'b0000101000000100001 : color = 12'he73;
15'b0000101000000100010 : color = 12'he73;
15'b0000101000000100011 : color = 12'he73;
15'b0000101000000100100 : color = 12'he51;
15'b0000101000000100101 : color = 12'hf00;
15'b0000101000000100110 : color = 12'hf42;
15'b0000101000000100111 : color = 12'he73;
15'b0000101000000101000 : color = 12'he73;
15'b0000101000000101001 : color = 12'he73;
15'b0000101000000101010 : color = 12'hf30;
15'b0000101000000101011 : color = 12'hf01;
15'b0000101000000101100 : color = 12'hf73;
15'b0000101000000101101 : color = 12'he73;
15'b0000101000000101110 : color = 12'he73;
15'b0000101000000101111 : color = 12'he73;
15'b0000101000000110000 : color = 12'he73;
15'b0000101000000110001 : color = 12'he73;
15'b0000101000000110010 : color = 12'he73;
15'b0000101000000110011 : color = 12'he72;
15'b0000101000000110100 : color = 12'hf10;
15'b0000101000000110101 : color = 12'hf63;
15'b0000101000000110110 : color = 12'he73;
15'b0000101000000110111 : color = 12'he73;
15'b0000101000000111000 : color = 12'he73;
15'b0000101000000111001 : color = 12'he73;
15'b0000101000000111010 : color = 12'he73;
15'b0000101000000111011 : color = 12'he73;
15'b0000101000000111100 : color = 12'he73;
15'b0000101000000111101 : color = 12'he73;
15'b0000101000000111110 : color = 12'he73;
15'b0000101000000111111 : color = 12'he73;
15'b0000101000001000000 : color = 12'he73;
15'b0000101000001000001 : color = 12'he73;
15'b0000101000001000010 : color = 12'he73;
15'b0000101000001000011 : color = 12'he73;
15'b0000101000001000100 : color = 12'he73;
15'b0000101000001000101 : color = 12'he73;
15'b0000101000001000110 : color = 12'he73;
15'b0000101000001000111 : color = 12'he73;
15'b0000101000001001000 : color = 12'he73;
15'b0000101000001001001 : color = 12'he73;
15'b0000101000001001010 : color = 12'he73;
15'b0000101000001001011 : color = 12'he73;
15'b0000101000001001100 : color = 12'he72;
15'b0000101000001001101 : color = 12'hf42;
15'b0000101000001001110 : color = 12'hf73;
15'b0000101000001001111 : color = 12'he73;
15'b0000101000001010000 : color = 12'he73;
15'b0000101000001010001 : color = 12'he61;
15'b0000101000001010010 : color = 12'hf00;
15'b0000101000001010011 : color = 12'hf53;
15'b0000101000001010100 : color = 12'he73;
15'b0000101000001010101 : color = 12'he73;
15'b0000101000001010110 : color = 12'he73;
15'b0000101000001010111 : color = 12'he73;
15'b0000101000001011000 : color = 12'he72;
15'b0000101000001011001 : color = 12'hf00;
15'b0000101000001011010 : color = 12'hf32;
15'b0000101000001011011 : color = 12'he73;
15'b0000101000001011100 : color = 12'he73;
15'b0000101000001011101 : color = 12'he73;
15'b0000101000001011110 : color = 12'he72;
15'b0000101000001011111 : color = 12'hf10;
15'b0000101000001100000 : color = 12'hf32;
15'b0000101000001100001 : color = 12'he73;
15'b0000101000001100010 : color = 12'he73;
15'b0000101000001100011 : color = 12'he73;
15'b0000101000001100100 : color = 12'he73;
15'b0000101000001100101 : color = 12'he73;
15'b0000101000001100110 : color = 12'he73;
15'b0000101000001100111 : color = 12'he73;
15'b0000101000001101000 : color = 12'he73;
15'b0000101000001101001 : color = 12'he73;
15'b0000101000001101010 : color = 12'he73;
15'b0000101000001101011 : color = 12'he73;
15'b0000101000001101100 : color = 12'he73;
15'b0000101000001101101 : color = 12'he73;
15'b0000101000001101110 : color = 12'he73;
15'b0000101000001101111 : color = 12'he73;
15'b0000101000001110000 : color = 12'he73;
15'b0000101000001110001 : color = 12'he73;
15'b0000101000001110010 : color = 12'he73;
15'b0000101000001110011 : color = 12'he73;
15'b0000101000001110100 : color = 12'he73;
15'b0000101000001110101 : color = 12'he73;
15'b0000101000001110110 : color = 12'he73;
15'b0000101000001110111 : color = 12'hf62;
15'b0000101000001111000 : color = 12'hf73;
15'b0000101000001111001 : color = 12'he73;
15'b0000101000001111010 : color = 12'he73;
15'b0000101000001111011 : color = 12'he73;
15'b0000101000001111100 : color = 12'he73;
15'b0000101000001111101 : color = 12'he73;
15'b0000101000001111110 : color = 12'he73;
15'b0000101000001111111 : color = 12'he73;
15'b0000101000010000000 : color = 12'he51;
15'b0000101000010000001 : color = 12'hf00;
15'b0000101000010000010 : color = 12'hf53;
15'b0000101000010000011 : color = 12'he73;
15'b0000101000010000100 : color = 12'he73;
15'b0000101000010000101 : color = 12'he73;
15'b0000101000010000110 : color = 12'he73;
15'b0000101000010000111 : color = 12'he73;
15'b0000101000010001000 : color = 12'he73;
15'b0000101000010001001 : color = 12'he73;
15'b0000101000010001010 : color = 12'he73;
15'b0000101000010001011 : color = 12'he73;
15'b0000101000010001100 : color = 12'he73;
15'b0000101000010001101 : color = 12'he73;
15'b0000101000010001110 : color = 12'he73;
15'b0000101000010001111 : color = 12'he73;
15'b0000101000010010000 : color = 12'he73;
15'b0000101000010010001 : color = 12'he73;
15'b0000101000010010010 : color = 12'he73;
15'b0000101000010010011 : color = 12'he73;
15'b0000101000010010100 : color = 12'he73;
15'b0000101000010010101 : color = 12'he73;
15'b0000101000010010110 : color = 12'he73;
15'b0000101000010010111 : color = 12'he73;
15'b0000101000010011000 : color = 12'he73;
15'b0000101000010011001 : color = 12'he73;
15'b0000101000010011010 : color = 12'he73;
15'b0000101000010011011 : color = 12'he73;
15'b0000101000010011100 : color = 12'he73;
15'b0000101000010011101 : color = 12'he73;
15'b0000101000010011110 : color = 12'he73;
15'b0000101000010011111 : color = 12'he73;
15'b0000101000010100000 : color = 12'he73;
15'b0000101000010100001 : color = 12'he73;
15'b0000101000010100010 : color = 12'he73;
15'b0000101000010100011 : color = 12'he73;
15'b0000101000010100100 : color = 12'he73;
15'b0000101000010100101 : color = 12'he73;
15'b0000101000010100110 : color = 12'he51;
15'b0000101000010100111 : color = 12'hf00;
15'b0000101000010101000 : color = 12'hf52;
15'b0000101000010101001 : color = 12'he73;
15'b0000101000010101010 : color = 12'he73;
15'b0000101000010101011 : color = 12'he73;
15'b0000101000010101100 : color = 12'he73;
15'b0000101000010101101 : color = 12'he73;
15'b0000101000010101110 : color = 12'he73;
15'b0000101000010101111 : color = 12'he73;
15'b0000101000010110000 : color = 12'he73;
15'b0000101000010110001 : color = 12'he72;
15'b0000101000010110010 : color = 12'hf00;
15'b0000101000010110011 : color = 12'hf00;
15'b0000101000010110100 : color = 12'hf63;
15'b0000101000010110101 : color = 12'he73;
15'b0000101000010110110 : color = 12'he73;
15'b0000101000010110111 : color = 12'hf40;
15'b0000101000010111000 : color = 12'hf01;
15'b0000101000010111001 : color = 12'hf73;
15'b0000101000010111010 : color = 12'he73;
15'b0000101000010111011 : color = 12'he73;
15'b0000101000010111100 : color = 12'he73;
15'b0000101000010111101 : color = 12'he73;
15'b0000101000010111110 : color = 12'he73;
15'b0000101000010111111 : color = 12'he73;
15'b0000101000011000000 : color = 12'he73;
15'b0000101000011000001 : color = 12'he73;
15'b0000101000011000010 : color = 12'he73;
15'b0000101000011000011 : color = 12'he73;
15'b0000101000011000100 : color = 12'he73;
15'b0000101000011000101 : color = 12'he73;
15'b0000101000011000110 : color = 12'he73;
15'b0000101000011000111 : color = 12'he73;
15'b0000101000011001000 : color = 12'he73;
15'b0000101000011001001 : color = 12'he73;
15'b0000101000011001010 : color = 12'he73;
15'b0000101000011001011 : color = 12'he73;
15'b0000101000011001100 : color = 12'he73;
15'b0000101000011001101 : color = 12'he62;
15'b0000101000011001110 : color = 12'hf63;
15'b0000101000011001111 : color = 12'he73;
15'b0000101000011010000 : color = 12'he73;
15'b0000101000011010001 : color = 12'he73;
15'b0000101000011010010 : color = 12'he73;
15'b0000101000011010011 : color = 12'he73;
15'b0000101000011010100 : color = 12'he73;
15'b0000101000011010101 : color = 12'he73;
15'b0000101000011010110 : color = 12'he73;
15'b0000101000011010111 : color = 12'he73;
15'b0000101000011011000 : color = 12'he73;
15'b0000101000011011001 : color = 12'he73;
15'b0000101000011011010 : color = 12'he73;
15'b0000101000011011011 : color = 12'he73;
15'b0000101000011011100 : color = 12'he73;
15'b0000101000011011101 : color = 12'he73;
15'b0000101000011011110 : color = 12'he73;
15'b0000101000011011111 : color = 12'he73;
15'b0000101000011100000 : color = 12'he73;
15'b0000101000011100001 : color = 12'he73;
15'b0000101000011100010 : color = 12'he73;
15'b0000101000011100011 : color = 12'he73;
15'b0000101000011100100 : color = 12'he73;
15'b0000101000011100101 : color = 12'he73;
15'b0000101000011100110 : color = 12'he73;
15'b0000101000011100111 : color = 12'he73;
15'b0000101000011101000 : color = 12'he73;
15'b0000101000011101001 : color = 12'he73;
15'b0000101000011101010 : color = 12'he73;
15'b0000101000011101011 : color = 12'he73;
15'b0000101000011101100 : color = 12'he73;
15'b0000101000011101101 : color = 12'he73;
15'b0000101000011101110 : color = 12'he73;
15'b0000101000011101111 : color = 12'he73;
15'b0000101000011110000 : color = 12'he73;
15'b0000101000011110001 : color = 12'he73;
15'b0000101000011110010 : color = 12'he73;
15'b0000101000011110011 : color = 12'he73;
15'b0000101000011110100 : color = 12'he73;
15'b0000101000011110101 : color = 12'he73;
15'b0000101000011110110 : color = 12'he73;
15'b0000101000011110111 : color = 12'he73;
15'b0000101000011111000 : color = 12'he73;
15'b0000101000011111001 : color = 12'he73;
15'b0000101000011111010 : color = 12'he73;
15'b0000101000011111011 : color = 12'he73;
15'b0000101000011111100 : color = 12'hf40;
15'b0000101000011111101 : color = 12'hf42;
15'b0000101000011111110 : color = 12'he73;
15'b0000101000011111111 : color = 12'he73;
15'b0000101000100000000 : color = 12'he73;
15'b0000101000100000001 : color = 12'hf41;
15'b0000101000100000010 : color = 12'hf63;
15'b0000101000100000011 : color = 12'he73;
15'b0000101000100000100 : color = 12'he73;
15'b0000101000100000101 : color = 12'he73;
15'b0000101000100000110 : color = 12'he73;
15'b0000101000100000111 : color = 12'he61;
15'b0000101000100001000 : color = 12'hf00;
15'b0000101000100001001 : color = 12'hf11;
15'b0000101000100001010 : color = 12'hf73;
15'b0000101000100001011 : color = 12'he73;
15'b0000101000100001100 : color = 12'he73;
15'b0000101000100001101 : color = 12'he73;
15'b0000101000100001110 : color = 12'he72;
15'b0000101000100001111 : color = 12'hf32;
15'b0000101000100010000 : color = 12'hf73;
15'b0000101000100010001 : color = 12'he73;
15'b0000101000100010010 : color = 12'he73;
15'b0000101000100010011 : color = 12'he73;
15'b0000101000100010100 : color = 12'he73;
15'b0000101000100010101 : color = 12'he73;
15'b0000101000100010110 : color = 12'he73;
15'b0000101000100010111 : color = 12'he73;
15'b0000101000100011000 : color = 12'he73;
15'b0000101000100011001 : color = 12'he73;
15'b0000101000100011010 : color = 12'he73;
15'b0000101000100011011 : color = 12'he73;
15'b0000101000100011100 : color = 12'he73;
15'b0000101000100011101 : color = 12'he73;
15'b0000101000100011110 : color = 12'he73;
15'b0000101000100011111 : color = 12'he73;
15'b0000101000100100000 : color = 12'he73;
15'b0000101000100100001 : color = 12'he73;
15'b0000101000100100010 : color = 12'he73;
15'b0000101000100100011 : color = 12'he73;
15'b0000101000100100100 : color = 12'he73;
15'b0000101000100100101 : color = 12'he73;
15'b0000101000100100110 : color = 12'he73;
15'b0000101000100100111 : color = 12'he73;
15'b0000101000100101000 : color = 12'he73;
15'b0000101000100101001 : color = 12'hf40;
15'b0000101000100101010 : color = 12'hf01;
15'b0000101000100101011 : color = 12'hf73;
15'b0000101000100101100 : color = 12'he73;
15'b0000101000100101101 : color = 12'hf40;
15'b0000101000100101110 : color = 12'hf32;
15'b0000101000100101111 : color = 12'hf73;
15'b0000101000100110000 : color = 12'he73;
15'b0000101000100110001 : color = 12'he73;
15'b0000101000100110010 : color = 12'he73;
15'b0000101000100110011 : color = 12'he73;
15'b0000101000100110100 : color = 12'he73;
15'b0000101000100110101 : color = 12'he51;
15'b0000101000100110110 : color = 12'hf00;
15'b0000101000100110111 : color = 12'hf53;
15'b0000101000100111000 : color = 12'he73;
15'b0000101000100111001 : color = 12'he73;
15'b0000101000100111010 : color = 12'he73;
15'b0000101000100111011 : color = 12'he73;
15'b0000101000100111100 : color = 12'he73;
15'b0000101000100111101 : color = 12'he73;
15'b0000101000100111110 : color = 12'he73;
15'b0000101000100111111 : color = 12'he73;
15'b0000101000101000000 : color = 12'he73;
15'b0000101000101000001 : color = 12'he73;
15'b0000101000101000010 : color = 12'he73;
15'b0000101000101000011 : color = 12'he73;
15'b0000101000101000100 : color = 12'he73;
15'b0000101000101000101 : color = 12'he73;
15'b0000101000101000110 : color = 12'he73;
15'b0000101000101000111 : color = 12'he73;
15'b0000101000101001000 : color = 12'he73;
15'b0000101000101001001 : color = 12'he73;
15'b0000101000101001010 : color = 12'he73;
15'b0000101000101001011 : color = 12'he73;
15'b0000101000101001100 : color = 12'he73;
15'b0000101000101001101 : color = 12'he73;
15'b0000101000101001110 : color = 12'he73;
15'b0000101000101001111 : color = 12'he73;
15'b0000101000101010000 : color = 12'he73;
15'b0000101000101010001 : color = 12'he72;
15'b0000101000101010010 : color = 12'hf31;
15'b0000101000101010011 : color = 12'hf73;
15'b0000101000101010100 : color = 12'he73;
15'b0000101000101010101 : color = 12'he73;
15'b0000101000101010110 : color = 12'he73;
15'b0000101000101010111 : color = 12'he61;
15'b0000101000101011000 : color = 12'hf00;
15'b0000101000101011001 : color = 12'hf53;
15'b0000101000101011010 : color = 12'he73;
15'b0000101000101011011 : color = 12'he61;
15'b0000101000101011100 : color = 12'hf11;
15'b0000101000101011101 : color = 12'hf63;
15'b0000101000101011110 : color = 12'he73;
15'b0000101000101011111 : color = 12'he73;
15'b0000101000101100000 : color = 12'he73;
15'b0000101000101100001 : color = 12'he73;
15'b0000101000101100010 : color = 12'he73;
15'b0000101000101100011 : color = 12'he51;
15'b0000101000101100100 : color = 12'hf00;
15'b0000101000101100101 : color = 12'hf53;
15'b0000101000101100110 : color = 12'he73;
15'b0000101000101100111 : color = 12'he73;
15'b0000101000101101000 : color = 12'he73;
15'b0000101000101101001 : color = 12'he73;
15'b0000101000101101010 : color = 12'he73;
15'b0000101000101101011 : color = 12'he73;
15'b0000101000101101100 : color = 12'he73;
15'b0000101000101101101 : color = 12'he73;
15'b0000101000101101110 : color = 12'he73;
15'b0000101000101101111 : color = 12'he73;
15'b0000101000101110000 : color = 12'he73;
15'b0000101000101110001 : color = 12'he73;
15'b0000101000101110010 : color = 12'he73;
15'b0000101000101110011 : color = 12'he73;
15'b0000101000101110100 : color = 12'he73;
15'b0000101000101110101 : color = 12'he73;
15'b0000101000101110110 : color = 12'he73;
15'b0000101000101110111 : color = 12'he73;
15'b0000101000101111000 : color = 12'he73;
15'b0000101000101111001 : color = 12'he73;
15'b0000101000101111010 : color = 12'he73;
15'b0000101000101111011 : color = 12'he73;
15'b0000101000101111100 : color = 12'he73;
15'b0000101000101111101 : color = 12'he73;
15'b0000101000101111110 : color = 12'he73;
15'b0000101000101111111 : color = 12'he73;
15'b0000101000110000000 : color = 12'he72;
15'b0000101000110000001 : color = 12'hf10;
15'b0000101000110000010 : color = 12'hf32;
15'b0000101000110000011 : color = 12'he73;
15'b0000101000110000100 : color = 12'he73;
15'b0000101000110000101 : color = 12'he73;
15'b0000101000110000110 : color = 12'he73;
15'b0000101000110000111 : color = 12'he61;
15'b0000101000110001000 : color = 12'hf00;
15'b0000101000110001001 : color = 12'hf63;
15'b0000101000110001010 : color = 12'he73;
15'b0000101000110001011 : color = 12'he73;
15'b0000101000110001100 : color = 12'he73;
15'b0000101000110001101 : color = 12'hf30;
15'b0000101000110001110 : color = 12'hf32;
15'b0000101000110001111 : color = 12'he73;
15'b0000101000110010000 : color = 12'he73;
15'b0000101000110010001 : color = 12'he73;
15'b0000101000110010010 : color = 12'he61;
15'b0000101000110010011 : color = 12'hf00;
15'b0000101000110010100 : color = 12'hf63;
15'b0000101000110010101 : color = 12'he73;
15'b0000101000110010110 : color = 12'he73;
15'b0000101000110010111 : color = 12'he73;
15'b0000101000110011000 : color = 12'he73;
15'b0000101000110011001 : color = 12'he73;
15'b0000101000110011010 : color = 12'he73;
15'b0000101000110011011 : color = 12'he73;
15'b0000101000110011100 : color = 12'he73;
15'b0000101000110011101 : color = 12'he73;
15'b0000101000110011110 : color = 12'he73;
15'b0000101000110011111 : color = 12'he73;
15'b0000101000110100000 : color = 12'he73;
15'b0000101000110100001 : color = 12'he73;
15'b0000101000110100010 : color = 12'he73;
15'b0000101000110100011 : color = 12'he73;
15'b0000101000110100100 : color = 12'he73;
15'b0000101000110100101 : color = 12'he73;
15'b0000101000110100110 : color = 12'he73;
15'b0000101000110100111 : color = 12'he73;
15'b0000101000110101000 : color = 12'he73;
15'b0000101000110101001 : color = 12'he73;
15'b0000101000110101010 : color = 12'he73;
15'b0000101000110101011 : color = 12'he73;
15'b0000101000110101100 : color = 12'he73;
15'b0000101000110101101 : color = 12'he73;
15'b0000101000110101110 : color = 12'he73;
15'b0000101000110101111 : color = 12'he73;
15'b0000101000110110000 : color = 12'he73;
15'b0000101000110110001 : color = 12'he62;
15'b0000101000110110010 : color = 12'hf10;
15'b0000101000110110011 : color = 12'hf11;
15'b0000101000110110100 : color = 12'hf73;
15'b0000101000110110101 : color = 12'he73;
15'b0000101000110110110 : color = 12'he73;
15'b0000101000110110111 : color = 12'he73;
15'b0000101000110111000 : color = 12'he73;
15'b0000101000110111001 : color = 12'he73;
15'b0000101000110111010 : color = 12'he73;
15'b0000101000110111011 : color = 12'hf40;
15'b0000101000110111100 : color = 12'hf32;
15'b0000101000110111101 : color = 12'hf73;
15'b0000101000110111110 : color = 12'he73;
15'b0000101000110111111 : color = 12'he73;
15'b0000101000111000000 : color = 12'he73;
15'b0000101000111000001 : color = 12'he73;
15'b0000101000111000010 : color = 12'he73;
15'b0000101000111000011 : color = 12'he73;
15'b0000101000111000100 : color = 12'he73;
15'b0000101000111000101 : color = 12'he73;
15'b0000101000111000110 : color = 12'he73;
15'b0000101000111000111 : color = 12'he73;
15'b0000101000111001000 : color = 12'he73;
15'b0000101000111001001 : color = 12'he73;
15'b0000101000111001010 : color = 12'he73;
15'b0000101000111001011 : color = 12'he73;
15'b0000101000111001100 : color = 12'he73;
15'b0000101000111001101 : color = 12'he73;
15'b0000101000111001110 : color = 12'he73;
15'b0000101000111001111 : color = 12'he73;
15'b0000101000111010000 : color = 12'he73;
15'b0000101000111010001 : color = 12'he73;
15'b0000101000111010010 : color = 12'he73;
15'b0000101000111010011 : color = 12'he73;
15'b0000101000111010100 : color = 12'he73;
15'b0000101000111010101 : color = 12'he73;
15'b0000101000111010110 : color = 12'he73;
15'b0000101000111010111 : color = 12'hf40;
15'b0000101000111011000 : color = 12'hf11;
15'b0000101000111011001 : color = 12'hf73;
15'b0000101000111011010 : color = 12'he73;
15'b0000101000111011011 : color = 12'he73;
15'b0000101000111011100 : color = 12'he72;
15'b0000101000111011101 : color = 12'hf00;
15'b0000101000111011110 : color = 12'hf32;
15'b0000101000111011111 : color = 12'hf73;
15'b0000101000111100000 : color = 12'he73;
15'b0000101000111100001 : color = 12'he73;
15'b0000101000111100010 : color = 12'he73;
15'b0000101000111100011 : color = 12'he72;
15'b0000101000111100100 : color = 12'hf00;
15'b0000101000111100101 : color = 12'hf00;
15'b0000101000111100110 : color = 12'hf42;
15'b0000101000111100111 : color = 12'he73;
15'b0000101000111101000 : color = 12'he73;
15'b0000101000111101001 : color = 12'he73;
15'b0000101000111101010 : color = 12'he73;
15'b0000101000111101011 : color = 12'he73;
15'b0000101000111101100 : color = 12'he73;
15'b0000101000111101101 : color = 12'he73;
15'b0000101000111101110 : color = 12'he73;
15'b0000101000111101111 : color = 12'he73;
15'b0000101000111110000 : color = 12'he73;
15'b0000101000111110001 : color = 12'he73;
15'b0000101000111110010 : color = 12'he73;
15'b0000101000111110011 : color = 12'he73;
15'b0000101000111110100 : color = 12'he73;
15'b0000101000111110101 : color = 12'he73;
15'b0000101000111110110 : color = 12'he73;
15'b0000101000111110111 : color = 12'he73;
15'b0000101000111111000 : color = 12'he73;
15'b0000101000111111001 : color = 12'he73;
15'b0000101000111111010 : color = 12'he73;
15'b0000101000111111011 : color = 12'he73;
15'b0000101000111111100 : color = 12'he73;
15'b0000101000111111101 : color = 12'he73;
15'b0000101000111111110 : color = 12'he73;
15'b0000101000000111101 : color = 12'he73;
15'b0000101000000111110 : color = 12'he73;
15'b0000101000000111111 : color = 12'he73;
15'b0000101000001000000 : color = 12'he73;
15'b0000101000001000001 : color = 12'he73;
15'b0000101000001000010 : color = 12'he73;
15'b0000101000001000011 : color = 12'he73;
15'b0000101000001000100 : color = 12'he73;
15'b0000101000001000101 : color = 12'he73;
15'b0000101000001000110 : color = 12'hf51;
15'b0000101000001000111 : color = 12'hf73;
15'b0000101000001001000 : color = 12'he73;
15'b0000101000001001001 : color = 12'he73;
15'b0000101000001001010 : color = 12'he73;
15'b0000101000001001011 : color = 12'he73;
15'b0000101000001001100 : color = 12'he73;
15'b0000101000001001101 : color = 12'hf40;
15'b0000101000001001110 : color = 12'hf00;
15'b0000101000001001111 : color = 12'hf63;
15'b0000101000001010000 : color = 12'he73;
15'b0000101000001010001 : color = 12'he73;
15'b0000101000001010010 : color = 12'he72;
15'b0000101000001010011 : color = 12'hf10;
15'b0000101000001010100 : color = 12'hf10;
15'b0000101000001010101 : color = 12'hf31;
15'b0000101000001010110 : color = 12'hf31;
15'b0000101000001010111 : color = 12'hf31;
15'b0000101000001011000 : color = 12'hf31;
15'b0000101000001011001 : color = 12'hf31;
15'b0000101000001011010 : color = 12'hf31;
15'b0000101000001011011 : color = 12'hf31;
15'b0000101000001011100 : color = 12'hf10;
15'b0000101000001011101 : color = 12'hf00;
15'b0000101000001011110 : color = 12'hf01;
15'b0000101000001011111 : color = 12'hf73;
15'b0000101000001100000 : color = 12'he73;
15'b0000101000001100001 : color = 12'he73;
15'b0000101000001100010 : color = 12'he73;
15'b0000101000001100011 : color = 12'he73;
15'b0000101000001100100 : color = 12'he73;
15'b0000101000001100101 : color = 12'he73;
15'b0000101000001100110 : color = 12'he73;
15'b0000101000001100111 : color = 12'he73;
15'b0000101000001101000 : color = 12'he73;
15'b0000101000001101001 : color = 12'he73;
15'b0000101000001101010 : color = 12'he73;
15'b0000101000001101011 : color = 12'he73;
15'b0000101000001101100 : color = 12'he73;
15'b0000101000001101101 : color = 12'he73;
15'b0000101000001101110 : color = 12'he73;
15'b0000101000001101111 : color = 12'he73;
15'b0000101000001110000 : color = 12'he73;
15'b0000101000001110001 : color = 12'he73;
15'b0000101000001110010 : color = 12'he73;
15'b0000101000001110011 : color = 12'he73;
15'b0000101000001110100 : color = 12'he73;
15'b0000101000001110101 : color = 12'he73;
15'b0000101000001110110 : color = 12'he73;
15'b0000101000001110111 : color = 12'he73;
15'b0000101000001111000 : color = 12'he73;
15'b0000101000001111001 : color = 12'he73;
15'b0000101000001111010 : color = 12'he61;
15'b0000101000001111011 : color = 12'hf00;
15'b0000101000001111100 : color = 12'hf53;
15'b0000101000001111101 : color = 12'he73;
15'b0000101000001111110 : color = 12'he73;
15'b0000101000001111111 : color = 12'he73;
15'b0000101000010000000 : color = 12'he73;
15'b0000101000010000001 : color = 12'he72;
15'b0000101000010000010 : color = 12'hf10;
15'b0000101000010000011 : color = 12'hf32;
15'b0000101000010000100 : color = 12'he73;
15'b0000101000010000101 : color = 12'he73;
15'b0000101000010000110 : color = 12'he73;
15'b0000101000010000111 : color = 12'he72;
15'b0000101000010001000 : color = 12'hf10;
15'b0000101000010001001 : color = 12'hf32;
15'b0000101000010001010 : color = 12'he73;
15'b0000101000010001011 : color = 12'he73;
15'b0000101000010001100 : color = 12'he73;
15'b0000101000010001101 : color = 12'he73;
15'b0000101000010001110 : color = 12'he73;
15'b0000101000010001111 : color = 12'he73;
15'b0000101000010010000 : color = 12'he73;
15'b0000101000010010001 : color = 12'he73;
15'b0000101000010010010 : color = 12'he73;
15'b0000101000010010011 : color = 12'he73;
15'b0000101000010010100 : color = 12'he73;
15'b0000101000010010101 : color = 12'he73;
15'b0000101000010010110 : color = 12'he73;
15'b0000101000010010111 : color = 12'he73;
15'b0000101000010011000 : color = 12'he73;
15'b0000101000010011001 : color = 12'he73;
15'b0000101000010011010 : color = 12'he73;
15'b0000101000010011011 : color = 12'he73;
15'b0000101000010011100 : color = 12'he73;
15'b0000101000010011101 : color = 12'he73;
15'b0000101000010011110 : color = 12'he73;
15'b0000101000010011111 : color = 12'he73;
15'b0000101000010100000 : color = 12'he73;
15'b0000101000010100001 : color = 12'he73;
15'b0000101000010100010 : color = 12'hf30;
15'b0000101000010100011 : color = 12'hf42;
15'b0000101000010100100 : color = 12'hf73;
15'b0000101000010100101 : color = 12'he73;
15'b0000101000010100110 : color = 12'he73;
15'b0000101000010100111 : color = 12'he73;
15'b0000101000010101000 : color = 12'he73;
15'b0000101000010101001 : color = 12'he51;
15'b0000101000010101010 : color = 12'hf00;
15'b0000101000010101011 : color = 12'hf53;
15'b0000101000010101100 : color = 12'he73;
15'b0000101000010101101 : color = 12'he73;
15'b0000101000010101110 : color = 12'he73;
15'b0000101000010101111 : color = 12'he73;
15'b0000101000010110000 : color = 12'he61;
15'b0000101000010110001 : color = 12'hf00;
15'b0000101000010110010 : color = 12'hf63;
15'b0000101000010110011 : color = 12'he73;
15'b0000101000010110100 : color = 12'he73;
15'b0000101000010110101 : color = 12'he73;
15'b0000101000010110110 : color = 12'he73;
15'b0000101000010110111 : color = 12'he73;
15'b0000101000010111000 : color = 12'he73;
15'b0000101000010111001 : color = 12'he73;
15'b0000101000010111010 : color = 12'he73;
15'b0000101000010111011 : color = 12'he73;
15'b0000101000010111100 : color = 12'he73;
15'b0000101000010111101 : color = 12'he73;
15'b0000101000010111110 : color = 12'he73;
15'b0000101000010111111 : color = 12'he73;
15'b0000101000011000000 : color = 12'he73;
15'b0000101000011000001 : color = 12'he73;
15'b0000101000011000010 : color = 12'he73;
15'b0000101000011000011 : color = 12'he73;
15'b0000101000011000100 : color = 12'he73;
15'b0000101000011000101 : color = 12'he73;
15'b0000101000011000110 : color = 12'he73;
15'b0000101000011000111 : color = 12'he73;
15'b0000101000011001000 : color = 12'he73;
15'b0000101000011001001 : color = 12'he73;
15'b0000101000011001010 : color = 12'he73;
15'b0000101000011001011 : color = 12'he73;
15'b0000101000011001100 : color = 12'he73;
15'b0000101000011001101 : color = 12'he73;
15'b0000101000011001110 : color = 12'he72;
15'b0000101000011001111 : color = 12'hf00;
15'b0000101000011010000 : color = 12'hf52;
15'b0000101000011010001 : color = 12'he73;
15'b0000101000011010010 : color = 12'he73;
15'b0000101000011010011 : color = 12'he72;
15'b0000101000011010100 : color = 12'hf31;
15'b0000101000011010101 : color = 12'hf63;
15'b0000101000011010110 : color = 12'he73;
15'b0000101000011010111 : color = 12'he73;
15'b0000101000011011000 : color = 12'he73;
15'b0000101000011011001 : color = 12'he73;
15'b0000101000011011010 : color = 12'he72;
15'b0000101000011011011 : color = 12'hf10;
15'b0000101000011011100 : color = 12'hf32;
15'b0000101000011011101 : color = 12'he73;
15'b0000101000011011110 : color = 12'he73;
15'b0000101000011011111 : color = 12'he73;
15'b0000101000011100000 : color = 12'hf40;
15'b0000101000011100001 : color = 12'hf01;
15'b0000101000011100010 : color = 12'hf73;
15'b0000101000011100011 : color = 12'he73;
15'b0000101000011100100 : color = 12'he73;
15'b0000101000011100101 : color = 12'he73;
15'b0000101000011100110 : color = 12'he73;
15'b0000101000011100111 : color = 12'he73;
15'b0000101000011101000 : color = 12'he73;
15'b0000101000011101001 : color = 12'he73;
15'b0000101000011101010 : color = 12'he73;
15'b0000101000011101011 : color = 12'he73;
15'b0000101000011101100 : color = 12'he73;
15'b0000101000011101101 : color = 12'he73;
15'b0000101000011101110 : color = 12'he73;
15'b0000101000011101111 : color = 12'he73;
15'b0000101000011110000 : color = 12'he73;
15'b0000101000011110001 : color = 12'he73;
15'b0000101000011110010 : color = 12'he73;
15'b0000101000011110011 : color = 12'he73;
15'b0000101000011110100 : color = 12'he73;
15'b0000101000011110101 : color = 12'he73;
15'b0000101000011110110 : color = 12'he73;
15'b0000101000011110111 : color = 12'he73;
15'b0000101000011111000 : color = 12'he73;
15'b0000101000011111001 : color = 12'he73;
15'b0000101000011111010 : color = 12'he73;
15'b0000101000011111011 : color = 12'he73;
15'b0000101000011111100 : color = 12'he73;
15'b0000101000011111101 : color = 12'hf30;
15'b0000101000011111110 : color = 12'hf32;
15'b0000101000011111111 : color = 12'hf73;
15'b0000101000100000000 : color = 12'he73;
15'b0000101000100000001 : color = 12'he73;
15'b0000101000100000010 : color = 12'he73;
15'b0000101000100000011 : color = 12'he73;
15'b0000101000100000100 : color = 12'he73;
15'b0000101000100000101 : color = 12'hf41;
15'b0000101000100000110 : color = 12'hf32;
15'b0000101000100000111 : color = 12'hf73;
15'b0000101000100001000 : color = 12'he73;
15'b0000101000100001001 : color = 12'he73;
15'b0000101000100001010 : color = 12'he73;
15'b0000101000100001011 : color = 12'he73;
15'b0000101000100001100 : color = 12'he73;
15'b0000101000100001101 : color = 12'he73;
15'b0000101000100001110 : color = 12'he73;
15'b0000101000100001111 : color = 12'he73;
15'b0000101000100010000 : color = 12'he73;
15'b0000101000100010001 : color = 12'he73;
15'b0000101000100010010 : color = 12'he73;
15'b0000101000100010011 : color = 12'he73;
15'b0000101000100010100 : color = 12'he73;
15'b0000101000100010101 : color = 12'he73;
15'b0000101000100010110 : color = 12'he73;
15'b0000101000100010111 : color = 12'he73;
15'b0000101000100011000 : color = 12'he73;
15'b0000101000100011001 : color = 12'he73;
15'b0000101000100011010 : color = 12'he73;
15'b0000101000100011011 : color = 12'he73;
15'b0000101000100011100 : color = 12'he73;
15'b0000101000100011101 : color = 12'he73;
15'b0000101000100011110 : color = 12'he73;
15'b0000101000100011111 : color = 12'he73;
15'b0000101000100100000 : color = 12'he73;
15'b0000101000100100001 : color = 12'he73;
15'b0000101000100100010 : color = 12'he73;
15'b0000101000100100011 : color = 12'he73;
15'b0000101000100100100 : color = 12'he73;
15'b0000101000100100101 : color = 12'he73;
15'b0000101000100100110 : color = 12'he73;
15'b0000101000100100111 : color = 12'he73;
15'b0000101000100101000 : color = 12'he73;
15'b0000101000100101001 : color = 12'he73;
15'b0000101000100101010 : color = 12'hf30;
15'b0000101000100101011 : color = 12'hf00;
15'b0000101000100101100 : color = 12'hf31;
15'b0000101000100101101 : color = 12'hf31;
15'b0000101000100101110 : color = 12'hf31;
15'b0000101000100101111 : color = 12'hf31;
15'b0000101000100110000 : color = 12'hf31;
15'b0000101000100110001 : color = 12'hf00;
15'b0000101000100110010 : color = 12'hf11;
15'b0000101000100110011 : color = 12'hf31;
15'b0000101000100110100 : color = 12'hf31;
15'b0000101000100110101 : color = 12'hf31;
15'b0000101000100110110 : color = 12'hf31;
15'b0000101000100110111 : color = 12'hf10;
15'b0000101000100111000 : color = 12'hf00;
15'b0000101000100111001 : color = 12'hf32;
15'b0000101000100111010 : color = 12'hf73;
15'b0000101000100111011 : color = 12'he73;
15'b0000101000100111100 : color = 12'he73;
15'b0000101000100111101 : color = 12'he73;
15'b0000101000100111110 : color = 12'he73;
15'b0000101000100111111 : color = 12'he73;
15'b0000101000101000000 : color = 12'he73;
15'b0000101000101000001 : color = 12'he73;
15'b0000101000101000010 : color = 12'he73;
15'b0000101000101000011 : color = 12'he73;
15'b0000101000101000100 : color = 12'he73;
15'b0000101000101000101 : color = 12'he73;
15'b0000101000101000110 : color = 12'he73;
15'b0000101000101000111 : color = 12'he73;
15'b0000101000101001000 : color = 12'he73;
15'b0000101000101001001 : color = 12'he73;
15'b0000101000101001010 : color = 12'he73;
15'b0000101000101001011 : color = 12'he73;
15'b0000101000101001100 : color = 12'he73;
15'b0000101000101001101 : color = 12'he73;
15'b0000101000101001110 : color = 12'he73;
15'b0000101000101001111 : color = 12'he73;
15'b0000101000101010000 : color = 12'he73;
15'b0000101000101010001 : color = 12'he73;
15'b0000101000101010010 : color = 12'hf40;
15'b0000101000101010011 : color = 12'hf01;
15'b0000101000101010100 : color = 12'hf73;
15'b0000101000101010101 : color = 12'he72;
15'b0000101000101010110 : color = 12'hf00;
15'b0000101000101010111 : color = 12'hf00;
15'b0000101000101011000 : color = 12'hf52;
15'b0000101000101011001 : color = 12'he73;
15'b0000101000101011010 : color = 12'he73;
15'b0000101000101011011 : color = 12'he73;
15'b0000101000101011100 : color = 12'he73;
15'b0000101000101011101 : color = 12'he73;
15'b0000101000101011110 : color = 12'he51;
15'b0000101000101011111 : color = 12'hf00;
15'b0000101000101100000 : color = 12'hf53;
15'b0000101000101100001 : color = 12'he73;
15'b0000101000101100010 : color = 12'he73;
15'b0000101000101100011 : color = 12'he73;
15'b0000101000101100100 : color = 12'he73;
15'b0000101000101100101 : color = 12'he73;
15'b0000101000101100110 : color = 12'he73;
15'b0000101000101100111 : color = 12'he73;
15'b0000101000101101000 : color = 12'he73;
15'b0000101000101101001 : color = 12'he73;
15'b0000101000101101010 : color = 12'he73;
15'b0000101000101101011 : color = 12'he73;
15'b0000101000101101100 : color = 12'he73;
15'b0000101000101101101 : color = 12'he73;
15'b0000101000101101110 : color = 12'he73;
15'b0000101000101101111 : color = 12'he73;
15'b0000101000101110000 : color = 12'he73;
15'b0000101000101110001 : color = 12'he73;
15'b0000101000101110010 : color = 12'he73;
15'b0000101000101110011 : color = 12'he73;
15'b0000101000101110100 : color = 12'he73;
15'b0000101000101110101 : color = 12'he73;
15'b0000101000101110110 : color = 12'he73;
15'b0000101000101110111 : color = 12'he73;
15'b0000101000101111000 : color = 12'he73;
15'b0000101000101111001 : color = 12'he72;
15'b0000101000101111010 : color = 12'hf42;
15'b0000101000101111011 : color = 12'hf73;
15'b0000101000101111100 : color = 12'he73;
15'b0000101000101111101 : color = 12'he73;
15'b0000101000101111110 : color = 12'he73;
15'b0000101000101111111 : color = 12'he73;
15'b0000101000110000000 : color = 12'he72;
15'b0000101000110000001 : color = 12'hf31;
15'b0000101000110000010 : color = 12'hf73;
15'b0000101000110000011 : color = 12'he73;
15'b0000101000110000100 : color = 12'he73;
15'b0000101000110000101 : color = 12'hf40;
15'b0000101000110000110 : color = 12'hf00;
15'b0000101000110000111 : color = 12'hf53;
15'b0000101000110001000 : color = 12'he73;
15'b0000101000110001001 : color = 12'he73;
15'b0000101000110001010 : color = 12'he73;
15'b0000101000110001011 : color = 12'he73;
15'b0000101000110001100 : color = 12'he72;
15'b0000101000110001101 : color = 12'hf31;
15'b0000101000110001110 : color = 12'hf73;
15'b0000101000110001111 : color = 12'he73;
15'b0000101000110010000 : color = 12'he73;
15'b0000101000110010001 : color = 12'he73;
15'b0000101000110010010 : color = 12'he73;
15'b0000101000110010011 : color = 12'he73;
15'b0000101000110010100 : color = 12'he73;
15'b0000101000110010101 : color = 12'he73;
15'b0000101000110010110 : color = 12'he73;
15'b0000101000110010111 : color = 12'he73;
15'b0000101000110011000 : color = 12'he73;
15'b0000101000110011001 : color = 12'he73;
15'b0000101000110011010 : color = 12'he73;
15'b0000101000110011011 : color = 12'he73;
15'b0000101000110011100 : color = 12'he73;
15'b0000101000110011101 : color = 12'he73;
15'b0000101000110011110 : color = 12'he73;
15'b0000101000110011111 : color = 12'he73;
15'b0000101000110100000 : color = 12'he73;
15'b0000101000110100001 : color = 12'he73;
15'b0000101000110100010 : color = 12'he73;
15'b0000101000110100011 : color = 12'he73;
15'b0000101000110100100 : color = 12'he73;
15'b0000101000110100101 : color = 12'he73;
15'b0000101000110100110 : color = 12'he73;
15'b0000101000110100111 : color = 12'he73;
15'b0000101000110101000 : color = 12'he73;
15'b0000101000110101001 : color = 12'he72;
15'b0000101000110101010 : color = 12'hf10;
15'b0000101000110101011 : color = 12'hf32;
15'b0000101000110101100 : color = 12'he73;
15'b0000101000110101101 : color = 12'he73;
15'b0000101000110101110 : color = 12'he73;
15'b0000101000110101111 : color = 12'he73;
15'b0000101000110110000 : color = 12'he61;
15'b0000101000110110001 : color = 12'hf00;
15'b0000101000110110010 : color = 12'hf63;
15'b0000101000110110011 : color = 12'he73;
15'b0000101000110110100 : color = 12'he73;
15'b0000101000110110101 : color = 12'he73;
15'b0000101000110110110 : color = 12'hf30;
15'b0000101000110110111 : color = 12'hf32;
15'b0000101000110111000 : color = 12'he73;
15'b0000101000110111001 : color = 12'he73;
15'b0000101000110111010 : color = 12'he73;
15'b0000101000110111011 : color = 12'he61;
15'b0000101000110111100 : color = 12'hf00;
15'b0000101000110111101 : color = 12'hf63;
15'b0000101000110111110 : color = 12'he73;
15'b0000101000110111111 : color = 12'he73;
15'b0000101000111000000 : color = 12'he73;
15'b0000101000111000001 : color = 12'he73;
15'b0000101000111000010 : color = 12'he73;
15'b0000101000111000011 : color = 12'he73;
15'b0000101000111000100 : color = 12'he73;
15'b0000101000111000101 : color = 12'he73;
15'b0000101000111000110 : color = 12'he73;
15'b0000101000111000111 : color = 12'he73;
15'b0000101000111001000 : color = 12'he73;
15'b0000101000111001001 : color = 12'he73;
15'b0000101000111001010 : color = 12'he73;
15'b0000101000111001011 : color = 12'he73;
15'b0000101000111001100 : color = 12'he73;
15'b0000101000111001101 : color = 12'he73;
15'b0000101000111001110 : color = 12'he73;
15'b0000101000111001111 : color = 12'he73;
15'b0000101000111010000 : color = 12'he73;
15'b0000101000111010001 : color = 12'he73;
15'b0000101000111010010 : color = 12'he73;
15'b0000101000111010011 : color = 12'he73;
15'b0000101000111010100 : color = 12'he73;
15'b0000101000111010101 : color = 12'he73;
15'b0000101000111010110 : color = 12'he73;
15'b0000101000111010111 : color = 12'he73;
15'b0000101000111011000 : color = 12'he73;
15'b0000101000111011001 : color = 12'hf51;
15'b0000101000111011010 : color = 12'hf00;
15'b0000101000111011011 : color = 12'hf42;
15'b0000101000111011100 : color = 12'he73;
15'b0000101000111011101 : color = 12'he73;
15'b0000101000111011110 : color = 12'he73;
15'b0000101000111011111 : color = 12'he73;
15'b0000101000111100000 : color = 12'he73;
15'b0000101000111100001 : color = 12'he73;
15'b0000101000111100010 : color = 12'he73;
15'b0000101000111100011 : color = 12'hf40;
15'b0000101000111100100 : color = 12'hf00;
15'b0000101000111100101 : color = 12'hf00;
15'b0000101000111100110 : color = 12'hf32;
15'b0000101000111100111 : color = 12'hf73;
15'b0000101000111101000 : color = 12'he73;
15'b0000101000111101001 : color = 12'he73;
15'b0000101000111101010 : color = 12'he73;
15'b0000101000111101011 : color = 12'he73;
15'b0000101000111101100 : color = 12'he73;
15'b0000101000111101101 : color = 12'he73;
15'b0000101000111101110 : color = 12'he73;
15'b0000101000111101111 : color = 12'he73;
15'b0000101000111110000 : color = 12'he73;
15'b0000101000111110001 : color = 12'he73;
15'b0000101000111110010 : color = 12'he73;
15'b0000101000111110011 : color = 12'he73;
15'b0000101000111110100 : color = 12'he73;
15'b0000101000111110101 : color = 12'he73;
15'b0000101000111110110 : color = 12'he73;
15'b0000101000111110111 : color = 12'he73;
15'b0000101000111111000 : color = 12'he73;
15'b0000101000111111001 : color = 12'he73;
15'b0000101000111111010 : color = 12'he73;
15'b0000101000111111011 : color = 12'he73;
15'b0000101000111111100 : color = 12'he73;
15'b0000101000111111101 : color = 12'he73;
15'b0000101000111111110 : color = 12'he73;
15'b0000101000111111111 : color = 12'he61;
15'b0000101001000000000 : color = 12'hf01;
15'b0000101001000000001 : color = 12'hf73;
15'b0000101001000000010 : color = 12'he73;
15'b0000101001000000011 : color = 12'he73;
15'b0000101001000000100 : color = 12'he73;
15'b0000101001000000101 : color = 12'hf40;
15'b0000101001000000110 : color = 12'hf00;
15'b0000101001000000111 : color = 12'hf11;
15'b0000101001000001000 : color = 12'hf63;
15'b0000101001000001001 : color = 12'he73;
15'b0000101001000001010 : color = 12'he73;
15'b0000101001000001011 : color = 12'he73;
15'b0000101001000001100 : color = 12'hf30;
15'b0000101001000001101 : color = 12'hf01;
15'b0000101001000001110 : color = 12'hf63;
15'b0000101001000001111 : color = 12'he73;
15'b0000101001000010000 : color = 12'he73;
15'b0000101001000010001 : color = 12'he73;
15'b0000101001000010010 : color = 12'he73;
15'b0000101001000010011 : color = 12'he73;
15'b0000101001000010100 : color = 12'he73;
15'b0000101001000010101 : color = 12'he73;
15'b0000101001000010110 : color = 12'he73;
15'b0000101001000010111 : color = 12'he73;
15'b0000101001000011000 : color = 12'he73;
15'b0000101001000011001 : color = 12'he73;
15'b0000101001000011010 : color = 12'he73;
15'b0000101001000011011 : color = 12'he73;
15'b0000101001000011100 : color = 12'he73;
15'b0000101001000011101 : color = 12'he73;
15'b0000101001000011110 : color = 12'he73;
15'b0000101001000011111 : color = 12'he73;
15'b0000101001000100000 : color = 12'he73;
15'b0000101001000100001 : color = 12'he73;
15'b0000101001000100010 : color = 12'he73;
15'b0000101001000100011 : color = 12'he73;
15'b0000101001000100100 : color = 12'he73;
15'b0000101001000100101 : color = 12'he73;
15'b0000101001000100110 : color = 12'he73;
15'b0000101001000100111 : color = 12'he73;
15'b0000101000001100110 : color = 12'he73;
15'b0000101000001100111 : color = 12'he73;
15'b0000101000001101000 : color = 12'he73;
15'b0000101000001101001 : color = 12'he73;
15'b0000101000001101010 : color = 12'he73;
15'b0000101000001101011 : color = 12'he73;
15'b0000101000001101100 : color = 12'he73;
15'b0000101000001101101 : color = 12'he73;
15'b0000101000001101110 : color = 12'he73;
15'b0000101000001101111 : color = 12'he72;
15'b0000101000001110000 : color = 12'hf31;
15'b0000101000001110001 : color = 12'hf73;
15'b0000101000001110010 : color = 12'he73;
15'b0000101000001110011 : color = 12'he73;
15'b0000101000001110100 : color = 12'he73;
15'b0000101000001110101 : color = 12'he72;
15'b0000101000001110110 : color = 12'hf10;
15'b0000101000001110111 : color = 12'hf11;
15'b0000101000001111000 : color = 12'hf73;
15'b0000101000001111001 : color = 12'he73;
15'b0000101000001111010 : color = 12'he73;
15'b0000101000001111011 : color = 12'he61;
15'b0000101000001111100 : color = 12'hf00;
15'b0000101000001111101 : color = 12'hf63;
15'b0000101000001111110 : color = 12'he72;
15'b0000101000001111111 : color = 12'hf42;
15'b0000101000010000000 : color = 12'hf73;
15'b0000101000010000001 : color = 12'he73;
15'b0000101000010000010 : color = 12'he73;
15'b0000101000010000011 : color = 12'he73;
15'b0000101000010000100 : color = 12'he73;
15'b0000101000010000101 : color = 12'hf30;
15'b0000101000010000110 : color = 12'hf00;
15'b0000101000010000111 : color = 12'hf42;
15'b0000101000010001000 : color = 12'hf73;
15'b0000101000010001001 : color = 12'he73;
15'b0000101000010001010 : color = 12'he73;
15'b0000101000010001011 : color = 12'he73;
15'b0000101000010001100 : color = 12'he73;
15'b0000101000010001101 : color = 12'he73;
15'b0000101000010001110 : color = 12'he73;
15'b0000101000010001111 : color = 12'he73;
15'b0000101000010010000 : color = 12'he73;
15'b0000101000010010001 : color = 12'he73;
15'b0000101000010010010 : color = 12'he73;
15'b0000101000010010011 : color = 12'he73;
15'b0000101000010010100 : color = 12'he73;
15'b0000101000010010101 : color = 12'he73;
15'b0000101000010010110 : color = 12'he73;
15'b0000101000010010111 : color = 12'he73;
15'b0000101000010011000 : color = 12'he73;
15'b0000101000010011001 : color = 12'he73;
15'b0000101000010011010 : color = 12'he73;
15'b0000101000010011011 : color = 12'he73;
15'b0000101000010011100 : color = 12'he73;
15'b0000101000010011101 : color = 12'he73;
15'b0000101000010011110 : color = 12'he73;
15'b0000101000010011111 : color = 12'he73;
15'b0000101000010100000 : color = 12'he73;
15'b0000101000010100001 : color = 12'he73;
15'b0000101000010100010 : color = 12'he73;
15'b0000101000010100011 : color = 12'he61;
15'b0000101000010100100 : color = 12'hf00;
15'b0000101000010100101 : color = 12'hf53;
15'b0000101000010100110 : color = 12'he73;
15'b0000101000010100111 : color = 12'he73;
15'b0000101000010101000 : color = 12'he73;
15'b0000101000010101001 : color = 12'he73;
15'b0000101000010101010 : color = 12'he72;
15'b0000101000010101011 : color = 12'hf10;
15'b0000101000010101100 : color = 12'hf32;
15'b0000101000010101101 : color = 12'he73;
15'b0000101000010101110 : color = 12'he73;
15'b0000101000010101111 : color = 12'he73;
15'b0000101000010110000 : color = 12'he72;
15'b0000101000010110001 : color = 12'hf10;
15'b0000101000010110010 : color = 12'hf32;
15'b0000101000010110011 : color = 12'he73;
15'b0000101000010110100 : color = 12'he73;
15'b0000101000010110101 : color = 12'he73;
15'b0000101000010110110 : color = 12'he73;
15'b0000101000010110111 : color = 12'he73;
15'b0000101000010111000 : color = 12'he73;
15'b0000101000010111001 : color = 12'he73;
15'b0000101000010111010 : color = 12'he73;
15'b0000101000010111011 : color = 12'he73;
15'b0000101000010111100 : color = 12'he73;
15'b0000101000010111101 : color = 12'he73;
15'b0000101000010111110 : color = 12'he73;
15'b0000101000010111111 : color = 12'he73;
15'b0000101000011000000 : color = 12'he73;
15'b0000101000011000001 : color = 12'he73;
15'b0000101000011000010 : color = 12'he73;
15'b0000101000011000011 : color = 12'he73;
15'b0000101000011000100 : color = 12'he73;
15'b0000101000011000101 : color = 12'he73;
15'b0000101000011000110 : color = 12'he73;
15'b0000101000011000111 : color = 12'he73;
15'b0000101000011001000 : color = 12'he73;
15'b0000101000011001001 : color = 12'he73;
15'b0000101000011001010 : color = 12'he73;
15'b0000101000011001011 : color = 12'he72;
15'b0000101000011001100 : color = 12'hf10;
15'b0000101000011001101 : color = 12'hf11;
15'b0000101000011001110 : color = 12'hf63;
15'b0000101000011001111 : color = 12'he73;
15'b0000101000011010000 : color = 12'he73;
15'b0000101000011010001 : color = 12'he73;
15'b0000101000011010010 : color = 12'he51;
15'b0000101000011010011 : color = 12'hf00;
15'b0000101000011010100 : color = 12'hf53;
15'b0000101000011010101 : color = 12'he73;
15'b0000101000011010110 : color = 12'he73;
15'b0000101000011010111 : color = 12'he73;
15'b0000101000011011000 : color = 12'he73;
15'b0000101000011011001 : color = 12'hf40;
15'b0000101000011011010 : color = 12'hf00;
15'b0000101000011011011 : color = 12'hf00;
15'b0000101000011011100 : color = 12'hf63;
15'b0000101000011011101 : color = 12'he73;
15'b0000101000011011110 : color = 12'he73;
15'b0000101000011011111 : color = 12'he73;
15'b0000101000011100000 : color = 12'he73;
15'b0000101000011100001 : color = 12'he73;
15'b0000101000011100010 : color = 12'he73;
15'b0000101000011100011 : color = 12'he73;
15'b0000101000011100100 : color = 12'he73;
15'b0000101000011100101 : color = 12'he73;
15'b0000101000011100110 : color = 12'he73;
15'b0000101000011100111 : color = 12'he73;
15'b0000101000011101000 : color = 12'he73;
15'b0000101000011101001 : color = 12'he73;
15'b0000101000011101010 : color = 12'he73;
15'b0000101000011101011 : color = 12'he73;
15'b0000101000011101100 : color = 12'he73;
15'b0000101000011101101 : color = 12'he73;
15'b0000101000011101110 : color = 12'he73;
15'b0000101000011101111 : color = 12'he73;
15'b0000101000011110000 : color = 12'he73;
15'b0000101000011110001 : color = 12'he73;
15'b0000101000011110010 : color = 12'he73;
15'b0000101000011110011 : color = 12'he73;
15'b0000101000011110100 : color = 12'he73;
15'b0000101000011110101 : color = 12'he73;
15'b0000101000011110110 : color = 12'he72;
15'b0000101000011110111 : color = 12'hf10;
15'b0000101000011111000 : color = 12'hf52;
15'b0000101000011111001 : color = 12'he73;
15'b0000101000011111010 : color = 12'he73;
15'b0000101000011111011 : color = 12'he73;
15'b0000101000011111100 : color = 12'he73;
15'b0000101000011111101 : color = 12'he72;
15'b0000101000011111110 : color = 12'hf00;
15'b0000101000011111111 : color = 12'hf42;
15'b0000101000100000000 : color = 12'he73;
15'b0000101000100000001 : color = 12'he73;
15'b0000101000100000010 : color = 12'he73;
15'b0000101000100000011 : color = 12'he72;
15'b0000101000100000100 : color = 12'hf10;
15'b0000101000100000101 : color = 12'hf32;
15'b0000101000100000110 : color = 12'he73;
15'b0000101000100000111 : color = 12'he73;
15'b0000101000100001000 : color = 12'he73;
15'b0000101000100001001 : color = 12'hf40;
15'b0000101000100001010 : color = 12'hf01;
15'b0000101000100001011 : color = 12'hf73;
15'b0000101000100001100 : color = 12'he73;
15'b0000101000100001101 : color = 12'he73;
15'b0000101000100001110 : color = 12'he73;
15'b0000101000100001111 : color = 12'he73;
15'b0000101000100010000 : color = 12'he73;
15'b0000101000100010001 : color = 12'he73;
15'b0000101000100010010 : color = 12'he73;
15'b0000101000100010011 : color = 12'he73;
15'b0000101000100010100 : color = 12'he73;
15'b0000101000100010101 : color = 12'he73;
15'b0000101000100010110 : color = 12'he73;
15'b0000101000100010111 : color = 12'he73;
15'b0000101000100011000 : color = 12'he73;
15'b0000101000100011001 : color = 12'he73;
15'b0000101000100011010 : color = 12'he73;
15'b0000101000100011011 : color = 12'he73;
15'b0000101000100011100 : color = 12'he73;
15'b0000101000100011101 : color = 12'he73;
15'b0000101000100011110 : color = 12'he73;
15'b0000101000100011111 : color = 12'he73;
15'b0000101000100100000 : color = 12'he73;
15'b0000101000100100001 : color = 12'he73;
15'b0000101000100100010 : color = 12'he73;
15'b0000101000100100011 : color = 12'he73;
15'b0000101000100100100 : color = 12'he73;
15'b0000101000100100101 : color = 12'hf40;
15'b0000101000100100110 : color = 12'hf00;
15'b0000101000100100111 : color = 12'hf00;
15'b0000101000100101000 : color = 12'hf42;
15'b0000101000100101001 : color = 12'he73;
15'b0000101000100101010 : color = 12'he73;
15'b0000101000100101011 : color = 12'he73;
15'b0000101000100101100 : color = 12'he73;
15'b0000101000100101101 : color = 12'he73;
15'b0000101000100101110 : color = 12'he73;
15'b0000101000100101111 : color = 12'hf51;
15'b0000101000100110000 : color = 12'hf00;
15'b0000101000100110001 : color = 12'hf32;
15'b0000101000100110010 : color = 12'hf73;
15'b0000101000100110011 : color = 12'he73;
15'b0000101000100110100 : color = 12'he73;
15'b0000101000100110101 : color = 12'he73;
15'b0000101000100110110 : color = 12'he73;
15'b0000101000100110111 : color = 12'he73;
15'b0000101000100111000 : color = 12'he73;
15'b0000101000100111001 : color = 12'he73;
15'b0000101000100111010 : color = 12'he73;
15'b0000101000100111011 : color = 12'he73;
15'b0000101000100111100 : color = 12'he73;
15'b0000101000100111101 : color = 12'he73;
15'b0000101000100111110 : color = 12'he73;
15'b0000101000100111111 : color = 12'he73;
15'b0000101000101000000 : color = 12'he73;
15'b0000101000101000001 : color = 12'he73;
15'b0000101000101000010 : color = 12'he73;
15'b0000101000101000011 : color = 12'he73;
15'b0000101000101000100 : color = 12'he73;
15'b0000101000101000101 : color = 12'he73;
15'b0000101000101000110 : color = 12'he73;
15'b0000101000101000111 : color = 12'he73;
15'b0000101000101001000 : color = 12'he73;
15'b0000101000101001001 : color = 12'he73;
15'b0000101000101001010 : color = 12'he73;
15'b0000101000101001011 : color = 12'he73;
15'b0000101000101001100 : color = 12'he73;
15'b0000101000101001101 : color = 12'he73;
15'b0000101000101001110 : color = 12'he73;
15'b0000101000101001111 : color = 12'he73;
15'b0000101000101010000 : color = 12'he73;
15'b0000101000101010001 : color = 12'he73;
15'b0000101000101010010 : color = 12'he73;
15'b0000101000101010011 : color = 12'hf30;
15'b0000101000101010100 : color = 12'hf11;
15'b0000101000101010101 : color = 12'hf73;
15'b0000101000101010110 : color = 12'he73;
15'b0000101000101010111 : color = 12'he73;
15'b0000101000101011000 : color = 12'he73;
15'b0000101000101011001 : color = 12'he61;
15'b0000101000101011010 : color = 12'hf00;
15'b0000101000101011011 : color = 12'hf53;
15'b0000101000101011100 : color = 12'he73;
15'b0000101000101011101 : color = 12'he73;
15'b0000101000101011110 : color = 12'he73;
15'b0000101000101011111 : color = 12'he73;
15'b0000101000101100000 : color = 12'he51;
15'b0000101000101100001 : color = 12'hf00;
15'b0000101000101100010 : color = 12'hf63;
15'b0000101000101100011 : color = 12'he73;
15'b0000101000101100100 : color = 12'he73;
15'b0000101000101100101 : color = 12'he73;
15'b0000101000101100110 : color = 12'he73;
15'b0000101000101100111 : color = 12'he73;
15'b0000101000101101000 : color = 12'he73;
15'b0000101000101101001 : color = 12'he73;
15'b0000101000101101010 : color = 12'he73;
15'b0000101000101101011 : color = 12'he73;
15'b0000101000101101100 : color = 12'he73;
15'b0000101000101101101 : color = 12'he73;
15'b0000101000101101110 : color = 12'he73;
15'b0000101000101101111 : color = 12'he73;
15'b0000101000101110000 : color = 12'he73;
15'b0000101000101110001 : color = 12'he73;
15'b0000101000101110010 : color = 12'he73;
15'b0000101000101110011 : color = 12'he73;
15'b0000101000101110100 : color = 12'he73;
15'b0000101000101110101 : color = 12'he73;
15'b0000101000101110110 : color = 12'he73;
15'b0000101000101110111 : color = 12'he73;
15'b0000101000101111000 : color = 12'hf41;
15'b0000101000101111001 : color = 12'hf73;
15'b0000101000101111010 : color = 12'he73;
15'b0000101000101111011 : color = 12'hf40;
15'b0000101000101111100 : color = 12'hf01;
15'b0000101000101111101 : color = 12'hf73;
15'b0000101000101111110 : color = 12'hf30;
15'b0000101000101111111 : color = 12'hf11;
15'b0000101000110000000 : color = 12'hf63;
15'b0000101000110000001 : color = 12'he73;
15'b0000101000110000010 : color = 12'he73;
15'b0000101000110000011 : color = 12'he73;
15'b0000101000110000100 : color = 12'he73;
15'b0000101000110000101 : color = 12'he73;
15'b0000101000110000110 : color = 12'he73;
15'b0000101000110000111 : color = 12'he51;
15'b0000101000110001000 : color = 12'hf00;
15'b0000101000110001001 : color = 12'hf53;
15'b0000101000110001010 : color = 12'he73;
15'b0000101000110001011 : color = 12'he73;
15'b0000101000110001100 : color = 12'he73;
15'b0000101000110001101 : color = 12'he73;
15'b0000101000110001110 : color = 12'he73;
15'b0000101000110001111 : color = 12'he73;
15'b0000101000110010000 : color = 12'he73;
15'b0000101000110010001 : color = 12'he73;
15'b0000101000110010010 : color = 12'he73;
15'b0000101000110010011 : color = 12'he73;
15'b0000101000110010100 : color = 12'he73;
15'b0000101000110010101 : color = 12'he73;
15'b0000101000110010110 : color = 12'he73;
15'b0000101000110010111 : color = 12'he73;
15'b0000101000110011000 : color = 12'he73;
15'b0000101000110011001 : color = 12'he73;
15'b0000101000110011010 : color = 12'he73;
15'b0000101000110011011 : color = 12'he73;
15'b0000101000110011100 : color = 12'he73;
15'b0000101000110011101 : color = 12'he73;
15'b0000101000110011110 : color = 12'he73;
15'b0000101000110011111 : color = 12'he73;
15'b0000101000110100000 : color = 12'he73;
15'b0000101000110100001 : color = 12'he73;
15'b0000101000110100010 : color = 12'he73;
15'b0000101000110100011 : color = 12'he73;
15'b0000101000110100100 : color = 12'he72;
15'b0000101000110100101 : color = 12'hf42;
15'b0000101000110100110 : color = 12'he73;
15'b0000101000110100111 : color = 12'he73;
15'b0000101000110101000 : color = 12'he73;
15'b0000101000110101001 : color = 12'he73;
15'b0000101000110101010 : color = 12'he73;
15'b0000101000110101011 : color = 12'he73;
15'b0000101000110101100 : color = 12'he73;
15'b0000101000110101101 : color = 12'he73;
15'b0000101000110101110 : color = 12'he61;
15'b0000101000110101111 : color = 12'hf00;
15'b0000101000110110000 : color = 12'hf42;
15'b0000101000110110001 : color = 12'he73;
15'b0000101000110110010 : color = 12'he73;
15'b0000101000110110011 : color = 12'he73;
15'b0000101000110110100 : color = 12'he73;
15'b0000101000110110101 : color = 12'he73;
15'b0000101000110110110 : color = 12'he73;
15'b0000101000110110111 : color = 12'he73;
15'b0000101000110111000 : color = 12'he73;
15'b0000101000110111001 : color = 12'he72;
15'b0000101000110111010 : color = 12'hf31;
15'b0000101000110111011 : color = 12'hf73;
15'b0000101000110111100 : color = 12'he73;
15'b0000101000110111101 : color = 12'he73;
15'b0000101000110111110 : color = 12'he73;
15'b0000101000110111111 : color = 12'he73;
15'b0000101000111000000 : color = 12'he73;
15'b0000101000111000001 : color = 12'he73;
15'b0000101000111000010 : color = 12'he73;
15'b0000101000111000011 : color = 12'he73;
15'b0000101000111000100 : color = 12'he73;
15'b0000101000111000101 : color = 12'he73;
15'b0000101000111000110 : color = 12'he73;
15'b0000101000111000111 : color = 12'he73;
15'b0000101000111001000 : color = 12'he73;
15'b0000101000111001001 : color = 12'he73;
15'b0000101000111001010 : color = 12'he73;
15'b0000101000111001011 : color = 12'he73;
15'b0000101000111001100 : color = 12'he73;
15'b0000101000111001101 : color = 12'he73;
15'b0000101000111001110 : color = 12'he73;
15'b0000101000111001111 : color = 12'he73;
15'b0000101000111010000 : color = 12'he73;
15'b0000101000111010001 : color = 12'he73;
15'b0000101000111010010 : color = 12'he72;
15'b0000101000111010011 : color = 12'hf10;
15'b0000101000111010100 : color = 12'hf32;
15'b0000101000111010101 : color = 12'he73;
15'b0000101000111010110 : color = 12'he73;
15'b0000101000111010111 : color = 12'he73;
15'b0000101000111011000 : color = 12'he73;
15'b0000101000111011001 : color = 12'he61;
15'b0000101000111011010 : color = 12'hf00;
15'b0000101000111011011 : color = 12'hf31;
15'b0000101000111011100 : color = 12'hf31;
15'b0000101000111011101 : color = 12'hf31;
15'b0000101000111011110 : color = 12'hf31;
15'b0000101000111011111 : color = 12'hf10;
15'b0000101000111100000 : color = 12'hf10;
15'b0000101000111100001 : color = 12'hf31;
15'b0000101000111100010 : color = 12'hf31;
15'b0000101000111100011 : color = 12'hf31;
15'b0000101000111100100 : color = 12'hf30;
15'b0000101000111100101 : color = 12'hf00;
15'b0000101000111100110 : color = 12'hf63;
15'b0000101000111100111 : color = 12'he73;
15'b0000101000111101000 : color = 12'he73;
15'b0000101000111101001 : color = 12'he73;
15'b0000101000111101010 : color = 12'he73;
15'b0000101000111101011 : color = 12'he73;
15'b0000101000111101100 : color = 12'he73;
15'b0000101000111101101 : color = 12'he73;
15'b0000101000111101110 : color = 12'he73;
15'b0000101000111101111 : color = 12'he73;
15'b0000101000111110000 : color = 12'he73;
15'b0000101000111110001 : color = 12'he73;
15'b0000101000111110010 : color = 12'he73;
15'b0000101000111110011 : color = 12'he73;
15'b0000101000111110100 : color = 12'he73;
15'b0000101000111110101 : color = 12'he73;
15'b0000101000111110110 : color = 12'he73;
15'b0000101000111110111 : color = 12'he73;
15'b0000101000111111000 : color = 12'he73;
15'b0000101000111111001 : color = 12'he73;
15'b0000101000111111010 : color = 12'he73;
15'b0000101000111111011 : color = 12'he73;
15'b0000101000111111100 : color = 12'he73;
15'b0000101000111111101 : color = 12'he73;
15'b0000101000111111110 : color = 12'he73;
15'b0000101000111111111 : color = 12'he73;
15'b0000101001000000000 : color = 12'he62;
15'b0000101001000000001 : color = 12'hf30;
15'b0000101001000000010 : color = 12'hf11;
15'b0000101001000000011 : color = 12'hf63;
15'b0000101001000000100 : color = 12'he73;
15'b0000101001000000101 : color = 12'he73;
15'b0000101001000000110 : color = 12'he73;
15'b0000101001000000111 : color = 12'he73;
15'b0000101001000001000 : color = 12'he73;
15'b0000101001000001001 : color = 12'he73;
15'b0000101001000001010 : color = 12'he72;
15'b0000101001000001011 : color = 12'hf30;
15'b0000101001000001100 : color = 12'hf00;
15'b0000101001000001101 : color = 12'hf31;
15'b0000101001000001110 : color = 12'hf63;
15'b0000101001000001111 : color = 12'he73;
15'b0000101001000010000 : color = 12'he73;
15'b0000101001000010001 : color = 12'he73;
15'b0000101001000010010 : color = 12'he73;
15'b0000101001000010011 : color = 12'he73;
15'b0000101001000010100 : color = 12'he73;
15'b0000101001000010101 : color = 12'he73;
15'b0000101001000010110 : color = 12'he73;
15'b0000101001000010111 : color = 12'he73;
15'b0000101001000011000 : color = 12'he73;
15'b0000101001000011001 : color = 12'he73;
15'b0000101001000011010 : color = 12'he73;
15'b0000101001000011011 : color = 12'he73;
15'b0000101001000011100 : color = 12'he73;
15'b0000101001000011101 : color = 12'he73;
15'b0000101001000011110 : color = 12'he73;
15'b0000101001000011111 : color = 12'he73;
15'b0000101001000100000 : color = 12'he73;
15'b0000101001000100001 : color = 12'he73;
15'b0000101001000100010 : color = 12'he73;
15'b0000101001000100011 : color = 12'he73;
15'b0000101001000100100 : color = 12'he73;
15'b0000101001000100101 : color = 12'he73;
15'b0000101001000100110 : color = 12'he73;
15'b0000101001000100111 : color = 12'he62;
15'b0000101001000101000 : color = 12'hf00;
15'b0000101001000101001 : color = 12'hf53;
15'b0000101001000101010 : color = 12'he73;
15'b0000101001000101011 : color = 12'he73;
15'b0000101001000101100 : color = 12'he73;
15'b0000101001000101101 : color = 12'he61;
15'b0000101001000101110 : color = 12'hf00;
15'b0000101001000101111 : color = 12'hf11;
15'b0000101001000110000 : color = 12'hf73;
15'b0000101001000110001 : color = 12'he73;
15'b0000101001000110010 : color = 12'he73;
15'b0000101001000110011 : color = 12'he73;
15'b0000101001000110100 : color = 12'he51;
15'b0000101001000110101 : color = 12'hf01;
15'b0000101001000110110 : color = 12'hf63;
15'b0000101001000110111 : color = 12'he73;
15'b0000101001000111000 : color = 12'he73;
15'b0000101001000111001 : color = 12'he61;
15'b0000101001000111010 : color = 12'hf42;
15'b0000101001000111011 : color = 12'hf73;
15'b0000101001000111100 : color = 12'he73;
15'b0000101001000111101 : color = 12'he73;
15'b0000101001000111110 : color = 12'he73;
15'b0000101001000111111 : color = 12'he73;
15'b0000101001001000000 : color = 12'he73;
15'b0000101001001000001 : color = 12'he73;
15'b0000101001001000010 : color = 12'he73;
15'b0000101001001000011 : color = 12'he73;
15'b0000101001001000100 : color = 12'he73;
15'b0000101001001000101 : color = 12'he73;
15'b0000101001001000110 : color = 12'he73;
15'b0000101001001000111 : color = 12'he73;
15'b0000101001001001000 : color = 12'he73;
15'b0000101001001001001 : color = 12'he73;
15'b0000101001001001010 : color = 12'he73;
15'b0000101001001001011 : color = 12'he73;
15'b0000101001001001100 : color = 12'he73;
15'b0000101001001001101 : color = 12'he73;
15'b0000101001001001110 : color = 12'he73;
15'b0000101001001001111 : color = 12'he73;
15'b0000101001001010000 : color = 12'he73;
15'b0000101000010001111 : color = 12'he73;
15'b0000101000010010000 : color = 12'he73;
15'b0000101000010010001 : color = 12'he73;
15'b0000101000010010010 : color = 12'he73;
15'b0000101000010010011 : color = 12'he73;
15'b0000101000010010100 : color = 12'he73;
15'b0000101000010010101 : color = 12'he73;
15'b0000101000010010110 : color = 12'he73;
15'b0000101000010010111 : color = 12'he73;
15'b0000101000010011000 : color = 12'he73;
15'b0000101000010011001 : color = 12'he72;
15'b0000101000010011010 : color = 12'hf11;
15'b0000101000010011011 : color = 12'hf73;
15'b0000101000010011100 : color = 12'he73;
15'b0000101000010011101 : color = 12'he73;
15'b0000101000010011110 : color = 12'he61;
15'b0000101000010011111 : color = 12'hf00;
15'b0000101000010100000 : color = 12'hf42;
15'b0000101000010100001 : color = 12'he73;
15'b0000101000010100010 : color = 12'he73;
15'b0000101000010100011 : color = 12'he73;
15'b0000101000010100100 : color = 12'hf40;
15'b0000101000010100101 : color = 12'hf32;
15'b0000101000010100110 : color = 12'he73;
15'b0000101000010100111 : color = 12'he72;
15'b0000101000010101000 : color = 12'hf10;
15'b0000101000010101001 : color = 12'hf00;
15'b0000101000010101010 : color = 12'hf52;
15'b0000101000010101011 : color = 12'he73;
15'b0000101000010101100 : color = 12'he73;
15'b0000101000010101101 : color = 12'he61;
15'b0000101000010101110 : color = 12'hf00;
15'b0000101000010101111 : color = 12'hf63;
15'b0000101000010110000 : color = 12'he73;
15'b0000101000010110001 : color = 12'he73;
15'b0000101000010110010 : color = 12'he73;
15'b0000101000010110011 : color = 12'he73;
15'b0000101000010110100 : color = 12'he73;
15'b0000101000010110101 : color = 12'he73;
15'b0000101000010110110 : color = 12'he73;
15'b0000101000010110111 : color = 12'he73;
15'b0000101000010111000 : color = 12'he73;
15'b0000101000010111001 : color = 12'he73;
15'b0000101000010111010 : color = 12'he73;
15'b0000101000010111011 : color = 12'he73;
15'b0000101000010111100 : color = 12'he73;
15'b0000101000010111101 : color = 12'he73;
15'b0000101000010111110 : color = 12'he73;
15'b0000101000010111111 : color = 12'he73;
15'b0000101000011000000 : color = 12'he73;
15'b0000101000011000001 : color = 12'he73;
15'b0000101000011000010 : color = 12'he73;
15'b0000101000011000011 : color = 12'he73;
15'b0000101000011000100 : color = 12'he73;
15'b0000101000011000101 : color = 12'he73;
15'b0000101000011000110 : color = 12'he73;
15'b0000101000011000111 : color = 12'he72;
15'b0000101000011001000 : color = 12'hf31;
15'b0000101000011001001 : color = 12'hf73;
15'b0000101000011001010 : color = 12'he73;
15'b0000101000011001011 : color = 12'he73;
15'b0000101000011001100 : color = 12'he61;
15'b0000101000011001101 : color = 12'hf00;
15'b0000101000011001110 : color = 12'hf53;
15'b0000101000011001111 : color = 12'he73;
15'b0000101000011010000 : color = 12'he73;
15'b0000101000011010001 : color = 12'he73;
15'b0000101000011010010 : color = 12'he73;
15'b0000101000011010011 : color = 12'he72;
15'b0000101000011010100 : color = 12'hf10;
15'b0000101000011010101 : color = 12'hf32;
15'b0000101000011010110 : color = 12'he73;
15'b0000101000011010111 : color = 12'he73;
15'b0000101000011011000 : color = 12'he73;
15'b0000101000011011001 : color = 12'he72;
15'b0000101000011011010 : color = 12'hf10;
15'b0000101000011011011 : color = 12'hf32;
15'b0000101000011011100 : color = 12'he73;
15'b0000101000011011101 : color = 12'he73;
15'b0000101000011011110 : color = 12'he73;
15'b0000101000011011111 : color = 12'he73;
15'b0000101000011100000 : color = 12'he73;
15'b0000101000011100001 : color = 12'he73;
15'b0000101000011100010 : color = 12'he73;
15'b0000101000011100011 : color = 12'he73;
15'b0000101000011100100 : color = 12'he73;
15'b0000101000011100101 : color = 12'he73;
15'b0000101000011100110 : color = 12'he73;
15'b0000101000011100111 : color = 12'he73;
15'b0000101000011101000 : color = 12'he73;
15'b0000101000011101001 : color = 12'he73;
15'b0000101000011101010 : color = 12'he73;
15'b0000101000011101011 : color = 12'he73;
15'b0000101000011101100 : color = 12'he73;
15'b0000101000011101101 : color = 12'he73;
15'b0000101000011101110 : color = 12'he73;
15'b0000101000011101111 : color = 12'he73;
15'b0000101000011110000 : color = 12'he73;
15'b0000101000011110001 : color = 12'he73;
15'b0000101000011110010 : color = 12'he73;
15'b0000101000011110011 : color = 12'he73;
15'b0000101000011110100 : color = 12'he73;
15'b0000101000011110101 : color = 12'he61;
15'b0000101000011110110 : color = 12'hf00;
15'b0000101000011110111 : color = 12'hf00;
15'b0000101000011111000 : color = 12'hf63;
15'b0000101000011111001 : color = 12'he73;
15'b0000101000011111010 : color = 12'he73;
15'b0000101000011111011 : color = 12'he51;
15'b0000101000011111100 : color = 12'hf00;
15'b0000101000011111101 : color = 12'hf53;
15'b0000101000011111110 : color = 12'he73;
15'b0000101000011111111 : color = 12'he73;
15'b0000101000100000000 : color = 12'he73;
15'b0000101000100000001 : color = 12'he61;
15'b0000101000100000010 : color = 12'hf00;
15'b0000101000100000011 : color = 12'hf11;
15'b0000101000100000100 : color = 12'hf73;
15'b0000101000100000101 : color = 12'he73;
15'b0000101000100000110 : color = 12'he73;
15'b0000101000100000111 : color = 12'he73;
15'b0000101000100001000 : color = 12'he73;
15'b0000101000100001001 : color = 12'he73;
15'b0000101000100001010 : color = 12'he73;
15'b0000101000100001011 : color = 12'he73;
15'b0000101000100001100 : color = 12'he73;
15'b0000101000100001101 : color = 12'he73;
15'b0000101000100001110 : color = 12'he73;
15'b0000101000100001111 : color = 12'he73;
15'b0000101000100010000 : color = 12'he73;
15'b0000101000100010001 : color = 12'he73;
15'b0000101000100010010 : color = 12'he73;
15'b0000101000100010011 : color = 12'he73;
15'b0000101000100010100 : color = 12'he73;
15'b0000101000100010101 : color = 12'he73;
15'b0000101000100010110 : color = 12'he73;
15'b0000101000100010111 : color = 12'he73;
15'b0000101000100011000 : color = 12'he73;
15'b0000101000100011001 : color = 12'he73;
15'b0000101000100011010 : color = 12'he73;
15'b0000101000100011011 : color = 12'he73;
15'b0000101000100011100 : color = 12'he73;
15'b0000101000100011101 : color = 12'he73;
15'b0000101000100011110 : color = 12'he62;
15'b0000101000100011111 : color = 12'hf10;
15'b0000101000100100000 : color = 12'hf53;
15'b0000101000100100001 : color = 12'he73;
15'b0000101000100100010 : color = 12'he73;
15'b0000101000100100011 : color = 12'he73;
15'b0000101000100100100 : color = 12'he73;
15'b0000101000100100101 : color = 12'he73;
15'b0000101000100100110 : color = 12'he73;
15'b0000101000100100111 : color = 12'he61;
15'b0000101000100101000 : color = 12'hf00;
15'b0000101000100101001 : color = 12'hf11;
15'b0000101000100101010 : color = 12'hf73;
15'b0000101000100101011 : color = 12'he73;
15'b0000101000100101100 : color = 12'he72;
15'b0000101000100101101 : color = 12'hf10;
15'b0000101000100101110 : color = 12'hf32;
15'b0000101000100101111 : color = 12'he73;
15'b0000101000100110000 : color = 12'he73;
15'b0000101000100110001 : color = 12'he73;
15'b0000101000100110010 : color = 12'hf40;
15'b0000101000100110011 : color = 12'hf01;
15'b0000101000100110100 : color = 12'hf73;
15'b0000101000100110101 : color = 12'he73;
15'b0000101000100110110 : color = 12'he73;
15'b0000101000100110111 : color = 12'he73;
15'b0000101000100111000 : color = 12'he73;
15'b0000101000100111001 : color = 12'he73;
15'b0000101000100111010 : color = 12'he73;
15'b0000101000100111011 : color = 12'he73;
15'b0000101000100111100 : color = 12'he73;
15'b0000101000100111101 : color = 12'he73;
15'b0000101000100111110 : color = 12'he73;
15'b0000101000100111111 : color = 12'he73;
15'b0000101000101000000 : color = 12'he73;
15'b0000101000101000001 : color = 12'he73;
15'b0000101000101000010 : color = 12'he73;
15'b0000101000101000011 : color = 12'he73;
15'b0000101000101000100 : color = 12'he73;
15'b0000101000101000101 : color = 12'he73;
15'b0000101000101000110 : color = 12'he73;
15'b0000101000101000111 : color = 12'he73;
15'b0000101000101001000 : color = 12'he73;
15'b0000101000101001001 : color = 12'he73;
15'b0000101000101001010 : color = 12'he73;
15'b0000101000101001011 : color = 12'he73;
15'b0000101000101001100 : color = 12'he73;
15'b0000101000101001101 : color = 12'he51;
15'b0000101000101001110 : color = 12'hf00;
15'b0000101000101001111 : color = 12'hf11;
15'b0000101000101010000 : color = 12'hf73;
15'b0000101000101010001 : color = 12'he73;
15'b0000101000101010010 : color = 12'he73;
15'b0000101000101010011 : color = 12'he73;
15'b0000101000101010100 : color = 12'he73;
15'b0000101000101010101 : color = 12'he73;
15'b0000101000101010110 : color = 12'he73;
15'b0000101000101010111 : color = 12'he73;
15'b0000101000101011000 : color = 12'he73;
15'b0000101000101011001 : color = 12'he62;
15'b0000101000101011010 : color = 12'hf10;
15'b0000101000101011011 : color = 12'hf00;
15'b0000101000101011100 : color = 12'hf42;
15'b0000101000101011101 : color = 12'he73;
15'b0000101000101011110 : color = 12'he73;
15'b0000101000101011111 : color = 12'he73;
15'b0000101000101100000 : color = 12'he73;
15'b0000101000101100001 : color = 12'he73;
15'b0000101000101100010 : color = 12'he73;
15'b0000101000101100011 : color = 12'he73;
15'b0000101000101100100 : color = 12'he73;
15'b0000101000101100101 : color = 12'he73;
15'b0000101000101100110 : color = 12'he73;
15'b0000101000101100111 : color = 12'he73;
15'b0000101000101101000 : color = 12'he73;
15'b0000101000101101001 : color = 12'he73;
15'b0000101000101101010 : color = 12'he73;
15'b0000101000101101011 : color = 12'he73;
15'b0000101000101101100 : color = 12'he73;
15'b0000101000101101101 : color = 12'he73;
15'b0000101000101101110 : color = 12'he73;
15'b0000101000101101111 : color = 12'he73;
15'b0000101000101110000 : color = 12'he73;
15'b0000101000101110001 : color = 12'he73;
15'b0000101000101110010 : color = 12'he73;
15'b0000101000101110011 : color = 12'he73;
15'b0000101000101110100 : color = 12'he73;
15'b0000101000101110101 : color = 12'he73;
15'b0000101000101110110 : color = 12'he73;
15'b0000101000101110111 : color = 12'he72;
15'b0000101000101111000 : color = 12'hf42;
15'b0000101000101111001 : color = 12'hf73;
15'b0000101000101111010 : color = 12'he73;
15'b0000101000101111011 : color = 12'he73;
15'b0000101000101111100 : color = 12'hf30;
15'b0000101000101111101 : color = 12'hf11;
15'b0000101000101111110 : color = 12'hf73;
15'b0000101000101111111 : color = 12'he73;
15'b0000101000110000000 : color = 12'he73;
15'b0000101000110000001 : color = 12'he73;
15'b0000101000110000010 : color = 12'he61;
15'b0000101000110000011 : color = 12'hf00;
15'b0000101000110000100 : color = 12'hf53;
15'b0000101000110000101 : color = 12'he73;
15'b0000101000110000110 : color = 12'he73;
15'b0000101000110000111 : color = 12'he73;
15'b0000101000110001000 : color = 12'he73;
15'b0000101000110001001 : color = 12'he51;
15'b0000101000110001010 : color = 12'hf00;
15'b0000101000110001011 : color = 12'hf63;
15'b0000101000110001100 : color = 12'he73;
15'b0000101000110001101 : color = 12'he73;
15'b0000101000110001110 : color = 12'he73;
15'b0000101000110001111 : color = 12'he73;
15'b0000101000110010000 : color = 12'he73;
15'b0000101000110010001 : color = 12'he73;
15'b0000101000110010010 : color = 12'he73;
15'b0000101000110010011 : color = 12'he73;
15'b0000101000110010100 : color = 12'he73;
15'b0000101000110010101 : color = 12'he73;
15'b0000101000110010110 : color = 12'he73;
15'b0000101000110010111 : color = 12'he73;
15'b0000101000110011000 : color = 12'he73;
15'b0000101000110011001 : color = 12'he73;
15'b0000101000110011010 : color = 12'he73;
15'b0000101000110011011 : color = 12'he73;
15'b0000101000110011100 : color = 12'he73;
15'b0000101000110011101 : color = 12'he73;
15'b0000101000110011110 : color = 12'he73;
15'b0000101000110011111 : color = 12'he73;
15'b0000101000110100000 : color = 12'he72;
15'b0000101000110100001 : color = 12'hf11;
15'b0000101000110100010 : color = 12'hf73;
15'b0000101000110100011 : color = 12'he73;
15'b0000101000110100100 : color = 12'hf40;
15'b0000101000110100101 : color = 12'hf01;
15'b0000101000110100110 : color = 12'hf40;
15'b0000101000110100111 : color = 12'hf32;
15'b0000101000110101000 : color = 12'hf73;
15'b0000101000110101001 : color = 12'he73;
15'b0000101000110101010 : color = 12'he73;
15'b0000101000110101011 : color = 12'he73;
15'b0000101000110101100 : color = 12'he73;
15'b0000101000110101101 : color = 12'he73;
15'b0000101000110101110 : color = 12'he73;
15'b0000101000110101111 : color = 12'he73;
15'b0000101000110110000 : color = 12'he51;
15'b0000101000110110001 : color = 12'hf00;
15'b0000101000110110010 : color = 12'hf53;
15'b0000101000110110011 : color = 12'he73;
15'b0000101000110110100 : color = 12'he73;
15'b0000101000110110101 : color = 12'he73;
15'b0000101000110110110 : color = 12'he73;
15'b0000101000110110111 : color = 12'he73;
15'b0000101000110111000 : color = 12'he73;
15'b0000101000110111001 : color = 12'he73;
15'b0000101000110111010 : color = 12'he73;
15'b0000101000110111011 : color = 12'he73;
15'b0000101000110111100 : color = 12'he73;
15'b0000101000110111101 : color = 12'he73;
15'b0000101000110111110 : color = 12'he73;
15'b0000101000110111111 : color = 12'he73;
15'b0000101000111000000 : color = 12'he73;
15'b0000101000111000001 : color = 12'he73;
15'b0000101000111000010 : color = 12'he73;
15'b0000101000111000011 : color = 12'he73;
15'b0000101000111000100 : color = 12'he73;
15'b0000101000111000101 : color = 12'he73;
15'b0000101000111000110 : color = 12'he73;
15'b0000101000111000111 : color = 12'he73;
15'b0000101000111001000 : color = 12'he73;
15'b0000101000111001001 : color = 12'he73;
15'b0000101000111001010 : color = 12'he73;
15'b0000101000111001011 : color = 12'he73;
15'b0000101000111001100 : color = 12'he73;
15'b0000101000111001101 : color = 12'he61;
15'b0000101000111001110 : color = 12'hf10;
15'b0000101000111001111 : color = 12'hf31;
15'b0000101000111010000 : color = 12'hf31;
15'b0000101000111010001 : color = 12'hf31;
15'b0000101000111010010 : color = 12'hf31;
15'b0000101000111010011 : color = 12'hf31;
15'b0000101000111010100 : color = 12'hf31;
15'b0000101000111010101 : color = 12'hf31;
15'b0000101000111010110 : color = 12'hf31;
15'b0000101000111010111 : color = 12'hf30;
15'b0000101000111011000 : color = 12'hf00;
15'b0000101000111011001 : color = 12'hf31;
15'b0000101000111011010 : color = 12'hf31;
15'b0000101000111011011 : color = 12'hf31;
15'b0000101000111011100 : color = 12'hf31;
15'b0000101000111011101 : color = 12'hf31;
15'b0000101000111011110 : color = 12'hf31;
15'b0000101000111011111 : color = 12'hf31;
15'b0000101000111100000 : color = 12'hf31;
15'b0000101000111100001 : color = 12'hf31;
15'b0000101000111100010 : color = 12'hf10;
15'b0000101000111100011 : color = 12'hf00;
15'b0000101000111100100 : color = 12'hf11;
15'b0000101000111100101 : color = 12'hf73;
15'b0000101000111100110 : color = 12'he73;
15'b0000101000111100111 : color = 12'he73;
15'b0000101000111101000 : color = 12'he73;
15'b0000101000111101001 : color = 12'he73;
15'b0000101000111101010 : color = 12'he73;
15'b0000101000111101011 : color = 12'he73;
15'b0000101000111101100 : color = 12'he73;
15'b0000101000111101101 : color = 12'he73;
15'b0000101000111101110 : color = 12'he73;
15'b0000101000111101111 : color = 12'he73;
15'b0000101000111110000 : color = 12'he73;
15'b0000101000111110001 : color = 12'he73;
15'b0000101000111110010 : color = 12'he73;
15'b0000101000111110011 : color = 12'he73;
15'b0000101000111110100 : color = 12'he73;
15'b0000101000111110101 : color = 12'he73;
15'b0000101000111110110 : color = 12'he73;
15'b0000101000111110111 : color = 12'he73;
15'b0000101000111111000 : color = 12'he73;
15'b0000101000111111001 : color = 12'he73;
15'b0000101000111111010 : color = 12'he73;
15'b0000101000111111011 : color = 12'he72;
15'b0000101000111111100 : color = 12'hf10;
15'b0000101000111111101 : color = 12'hf32;
15'b0000101000111111110 : color = 12'he73;
15'b0000101000111111111 : color = 12'he73;
15'b0000101001000000000 : color = 12'he73;
15'b0000101001000000001 : color = 12'he73;
15'b0000101001000000010 : color = 12'he61;
15'b0000101001000000011 : color = 12'hf00;
15'b0000101001000000100 : color = 12'hf63;
15'b0000101001000000101 : color = 12'he73;
15'b0000101001000000110 : color = 12'he73;
15'b0000101001000000111 : color = 12'he73;
15'b0000101001000001000 : color = 12'hf30;
15'b0000101001000001001 : color = 12'hf32;
15'b0000101001000001010 : color = 12'he73;
15'b0000101001000001011 : color = 12'he73;
15'b0000101001000001100 : color = 12'he73;
15'b0000101001000001101 : color = 12'he61;
15'b0000101001000001110 : color = 12'hf00;
15'b0000101001000001111 : color = 12'hf63;
15'b0000101001000010000 : color = 12'he73;
15'b0000101001000010001 : color = 12'he73;
15'b0000101001000010010 : color = 12'he73;
15'b0000101001000010011 : color = 12'he73;
15'b0000101001000010100 : color = 12'he73;
15'b0000101001000010101 : color = 12'he73;
15'b0000101001000010110 : color = 12'he73;
15'b0000101001000010111 : color = 12'he73;
15'b0000101001000011000 : color = 12'he73;
15'b0000101001000011001 : color = 12'he73;
15'b0000101001000011010 : color = 12'he73;
15'b0000101001000011011 : color = 12'he73;
15'b0000101001000011100 : color = 12'he73;
15'b0000101001000011101 : color = 12'he73;
15'b0000101001000011110 : color = 12'he73;
15'b0000101001000011111 : color = 12'he73;
15'b0000101001000100000 : color = 12'he73;
15'b0000101001000100001 : color = 12'he73;
15'b0000101001000100010 : color = 12'he73;
15'b0000101001000100011 : color = 12'he73;
15'b0000101001000100100 : color = 12'he73;
15'b0000101001000100101 : color = 12'he73;
15'b0000101001000100110 : color = 12'he73;
15'b0000101001000100111 : color = 12'he73;
15'b0000101001000101000 : color = 12'hf40;
15'b0000101001000101001 : color = 12'hf00;
15'b0000101001000101010 : color = 12'hf00;
15'b0000101001000101011 : color = 12'hf10;
15'b0000101001000101100 : color = 12'hf10;
15'b0000101001000101101 : color = 12'hf10;
15'b0000101001000101110 : color = 12'hf10;
15'b0000101001000101111 : color = 12'hf00;
15'b0000101001000110000 : color = 12'hf10;
15'b0000101001000110001 : color = 12'hf10;
15'b0000101001000110010 : color = 12'hf10;
15'b0000101001000110011 : color = 12'hf00;
15'b0000101001000110100 : color = 12'hf11;
15'b0000101001000110101 : color = 12'hf52;
15'b0000101001000110110 : color = 12'he73;
15'b0000101001000110111 : color = 12'he73;
15'b0000101001000111000 : color = 12'he73;
15'b0000101001000111001 : color = 12'he73;
15'b0000101001000111010 : color = 12'he73;
15'b0000101001000111011 : color = 12'he73;
15'b0000101001000111100 : color = 12'he73;
15'b0000101001000111101 : color = 12'he73;
15'b0000101001000111110 : color = 12'he73;
15'b0000101001000111111 : color = 12'he73;
15'b0000101001001000000 : color = 12'he73;
15'b0000101001001000001 : color = 12'he73;
15'b0000101001001000010 : color = 12'he73;
15'b0000101001001000011 : color = 12'he73;
15'b0000101001001000100 : color = 12'he73;
15'b0000101001001000101 : color = 12'he73;
15'b0000101001001000110 : color = 12'he73;
15'b0000101001001000111 : color = 12'he73;
15'b0000101001001001000 : color = 12'he73;
15'b0000101001001001001 : color = 12'he73;
15'b0000101001001001010 : color = 12'he73;
15'b0000101001001001011 : color = 12'he73;
15'b0000101001001001100 : color = 12'he73;
15'b0000101001001001101 : color = 12'he73;
15'b0000101001001001110 : color = 12'he73;
15'b0000101001001001111 : color = 12'he72;
15'b0000101001001010000 : color = 12'hf00;
15'b0000101001001010001 : color = 12'hf00;
15'b0000101001001010010 : color = 12'hf10;
15'b0000101001001010011 : color = 12'hf10;
15'b0000101001001010100 : color = 12'hf00;
15'b0000101001001010101 : color = 12'hf31;
15'b0000101001001010110 : color = 12'hf00;
15'b0000101001001010111 : color = 12'hf01;
15'b0000101001001011000 : color = 12'hf73;
15'b0000101001001011001 : color = 12'he73;
15'b0000101001001011010 : color = 12'he73;
15'b0000101001001011011 : color = 12'he73;
15'b0000101001001011100 : color = 12'he72;
15'b0000101001001011101 : color = 12'hf10;
15'b0000101001001011110 : color = 12'hf63;
15'b0000101001001011111 : color = 12'he73;
15'b0000101001001100000 : color = 12'he73;
15'b0000101001001100001 : color = 12'he73;
15'b0000101001001100010 : color = 12'he73;
15'b0000101001001100011 : color = 12'hf51;
15'b0000101001001100100 : color = 12'hf00;
15'b0000101001001100101 : color = 12'hf42;
15'b0000101001001100110 : color = 12'hf73;
15'b0000101001001100111 : color = 12'he73;
15'b0000101001001101000 : color = 12'he73;
15'b0000101001001101001 : color = 12'he73;
15'b0000101001001101010 : color = 12'he73;
15'b0000101001001101011 : color = 12'he73;
15'b0000101001001101100 : color = 12'he73;
15'b0000101001001101101 : color = 12'he73;
15'b0000101001001101110 : color = 12'he73;
15'b0000101001001101111 : color = 12'he73;
15'b0000101001001110000 : color = 12'he73;
15'b0000101001001110001 : color = 12'he73;
15'b0000101001001110010 : color = 12'he73;
15'b0000101001001110011 : color = 12'he73;
15'b0000101001001110100 : color = 12'he73;
15'b0000101001001110101 : color = 12'he73;
15'b0000101001001110110 : color = 12'he73;
15'b0000101001001110111 : color = 12'he73;
15'b0000101001001111000 : color = 12'he73;
15'b0000101001001111001 : color = 12'he73;
15'b0000101000010111000 : color = 12'he73;
15'b0000101000010111001 : color = 12'he73;
15'b0000101000010111010 : color = 12'he73;
15'b0000101000010111011 : color = 12'he73;
15'b0000101000010111100 : color = 12'he73;
15'b0000101000010111101 : color = 12'he73;
15'b0000101000010111110 : color = 12'he73;
15'b0000101000010111111 : color = 12'he73;
15'b0000101000011000000 : color = 12'he73;
15'b0000101000011000001 : color = 12'he73;
15'b0000101000011000010 : color = 12'he73;
15'b0000101000011000011 : color = 12'he51;
15'b0000101000011000100 : color = 12'hf11;
15'b0000101000011000101 : color = 12'hf73;
15'b0000101000011000110 : color = 12'he73;
15'b0000101000011000111 : color = 12'he51;
15'b0000101000011001000 : color = 12'hf00;
15'b0000101000011001001 : color = 12'hf63;
15'b0000101000011001010 : color = 12'he73;
15'b0000101000011001011 : color = 12'he73;
15'b0000101000011001100 : color = 12'he72;
15'b0000101000011001101 : color = 12'hf00;
15'b0000101000011001110 : color = 12'hf63;
15'b0000101000011001111 : color = 12'he73;
15'b0000101000011010000 : color = 12'he72;
15'b0000101000011010001 : color = 12'hf10;
15'b0000101000011010010 : color = 12'hf01;
15'b0000101000011010011 : color = 12'hf73;
15'b0000101000011010100 : color = 12'he73;
15'b0000101000011010101 : color = 12'he73;
15'b0000101000011010110 : color = 12'hf40;
15'b0000101000011010111 : color = 12'hf53;
15'b0000101000011011000 : color = 12'he73;
15'b0000101000011011001 : color = 12'he73;
15'b0000101000011011010 : color = 12'he73;
15'b0000101000011011011 : color = 12'he73;
15'b0000101000011011100 : color = 12'he73;
15'b0000101000011011101 : color = 12'he73;
15'b0000101000011011110 : color = 12'he73;
15'b0000101000011011111 : color = 12'he73;
15'b0000101000011100000 : color = 12'he73;
15'b0000101000011100001 : color = 12'he73;
15'b0000101000011100010 : color = 12'he73;
15'b0000101000011100011 : color = 12'he73;
15'b0000101000011100100 : color = 12'he73;
15'b0000101000011100101 : color = 12'he73;
15'b0000101000011100110 : color = 12'he73;
15'b0000101000011100111 : color = 12'he73;
15'b0000101000011101000 : color = 12'he73;
15'b0000101000011101001 : color = 12'he73;
15'b0000101000011101010 : color = 12'he73;
15'b0000101000011101011 : color = 12'he73;
15'b0000101000011101100 : color = 12'he61;
15'b0000101000011101101 : color = 12'hf31;
15'b0000101000011101110 : color = 12'hf31;
15'b0000101000011101111 : color = 12'hf31;
15'b0000101000011110000 : color = 12'hf10;
15'b0000101000011110001 : color = 12'hf00;
15'b0000101000011110010 : color = 12'hf11;
15'b0000101000011110011 : color = 12'hf73;
15'b0000101000011110100 : color = 12'he73;
15'b0000101000011110101 : color = 12'he61;
15'b0000101000011110110 : color = 12'hf00;
15'b0000101000011110111 : color = 12'hf53;
15'b0000101000011111000 : color = 12'he73;
15'b0000101000011111001 : color = 12'he73;
15'b0000101000011111010 : color = 12'he73;
15'b0000101000011111011 : color = 12'he73;
15'b0000101000011111100 : color = 12'he72;
15'b0000101000011111101 : color = 12'hf10;
15'b0000101000011111110 : color = 12'hf32;
15'b0000101000011111111 : color = 12'he73;
15'b0000101000100000000 : color = 12'he73;
15'b0000101000100000001 : color = 12'he73;
15'b0000101000100000010 : color = 12'he72;
15'b0000101000100000011 : color = 12'hf10;
15'b0000101000100000100 : color = 12'hf32;
15'b0000101000100000101 : color = 12'he73;
15'b0000101000100000110 : color = 12'he73;
15'b0000101000100000111 : color = 12'he73;
15'b0000101000100001000 : color = 12'he73;
15'b0000101000100001001 : color = 12'he73;
15'b0000101000100001010 : color = 12'he73;
15'b0000101000100001011 : color = 12'he73;
15'b0000101000100001100 : color = 12'he73;
15'b0000101000100001101 : color = 12'he73;
15'b0000101000100001110 : color = 12'he73;
15'b0000101000100001111 : color = 12'he73;
15'b0000101000100010000 : color = 12'he73;
15'b0000101000100010001 : color = 12'he73;
15'b0000101000100010010 : color = 12'he73;
15'b0000101000100010011 : color = 12'he73;
15'b0000101000100010100 : color = 12'he73;
15'b0000101000100010101 : color = 12'he73;
15'b0000101000100010110 : color = 12'he73;
15'b0000101000100010111 : color = 12'he73;
15'b0000101000100011000 : color = 12'he73;
15'b0000101000100011001 : color = 12'he73;
15'b0000101000100011010 : color = 12'he73;
15'b0000101000100011011 : color = 12'he73;
15'b0000101000100011100 : color = 12'he73;
15'b0000101000100011101 : color = 12'he73;
15'b0000101000100011110 : color = 12'he73;
15'b0000101000100011111 : color = 12'hf30;
15'b0000101000100100000 : color = 12'hf00;
15'b0000101000100100001 : color = 12'hf32;
15'b0000101000100100010 : color = 12'he73;
15'b0000101000100100011 : color = 12'he73;
15'b0000101000100100100 : color = 12'he51;
15'b0000101000100100101 : color = 12'hf00;
15'b0000101000100100110 : color = 12'hf53;
15'b0000101000100100111 : color = 12'he73;
15'b0000101000100101000 : color = 12'he73;
15'b0000101000100101001 : color = 12'he73;
15'b0000101000100101010 : color = 12'hf30;
15'b0000101000100101011 : color = 12'hf01;
15'b0000101000100101100 : color = 12'hf73;
15'b0000101000100101101 : color = 12'he73;
15'b0000101000100101110 : color = 12'he73;
15'b0000101000100101111 : color = 12'he73;
15'b0000101000100110000 : color = 12'he73;
15'b0000101000100110001 : color = 12'he73;
15'b0000101000100110010 : color = 12'he73;
15'b0000101000100110011 : color = 12'he73;
15'b0000101000100110100 : color = 12'he73;
15'b0000101000100110101 : color = 12'he73;
15'b0000101000100110110 : color = 12'he73;
15'b0000101000100110111 : color = 12'he73;
15'b0000101000100111000 : color = 12'he73;
15'b0000101000100111001 : color = 12'he73;
15'b0000101000100111010 : color = 12'he73;
15'b0000101000100111011 : color = 12'he73;
15'b0000101000100111100 : color = 12'he73;
15'b0000101000100111101 : color = 12'he73;
15'b0000101000100111110 : color = 12'he73;
15'b0000101000100111111 : color = 12'he73;
15'b0000101000101000000 : color = 12'he73;
15'b0000101000101000001 : color = 12'he73;
15'b0000101000101000010 : color = 12'he73;
15'b0000101000101000011 : color = 12'he73;
15'b0000101000101000100 : color = 12'he73;
15'b0000101000101000101 : color = 12'he72;
15'b0000101000101000110 : color = 12'hf30;
15'b0000101000101000111 : color = 12'hf00;
15'b0000101000101001000 : color = 12'hf11;
15'b0000101000101001001 : color = 12'hf31;
15'b0000101000101001010 : color = 12'hf31;
15'b0000101000101001011 : color = 12'hf31;
15'b0000101000101001100 : color = 12'hf31;
15'b0000101000101001101 : color = 12'hf30;
15'b0000101000101001110 : color = 12'hf10;
15'b0000101000101001111 : color = 12'hf10;
15'b0000101000101010000 : color = 12'hf10;
15'b0000101000101010001 : color = 12'hf00;
15'b0000101000101010010 : color = 12'hf00;
15'b0000101000101010011 : color = 12'hf11;
15'b0000101000101010100 : color = 12'hf73;
15'b0000101000101010101 : color = 12'he72;
15'b0000101000101010110 : color = 12'hf10;
15'b0000101000101010111 : color = 12'hf32;
15'b0000101000101011000 : color = 12'he73;
15'b0000101000101011001 : color = 12'he73;
15'b0000101000101011010 : color = 12'he73;
15'b0000101000101011011 : color = 12'hf40;
15'b0000101000101011100 : color = 12'hf01;
15'b0000101000101011101 : color = 12'hf73;
15'b0000101000101011110 : color = 12'he73;
15'b0000101000101011111 : color = 12'he73;
15'b0000101000101100000 : color = 12'he73;
15'b0000101000101100001 : color = 12'he73;
15'b0000101000101100010 : color = 12'he73;
15'b0000101000101100011 : color = 12'he73;
15'b0000101000101100100 : color = 12'he73;
15'b0000101000101100101 : color = 12'he73;
15'b0000101000101100110 : color = 12'he73;
15'b0000101000101100111 : color = 12'he73;
15'b0000101000101101000 : color = 12'he73;
15'b0000101000101101001 : color = 12'he73;
15'b0000101000101101010 : color = 12'he73;
15'b0000101000101101011 : color = 12'he73;
15'b0000101000101101100 : color = 12'he73;
15'b0000101000101101101 : color = 12'he73;
15'b0000101000101101110 : color = 12'he73;
15'b0000101000101101111 : color = 12'he73;
15'b0000101000101110000 : color = 12'he73;
15'b0000101000101110001 : color = 12'he73;
15'b0000101000101110010 : color = 12'he73;
15'b0000101000101110011 : color = 12'he73;
15'b0000101000101110100 : color = 12'he73;
15'b0000101000101110101 : color = 12'he61;
15'b0000101000101110110 : color = 12'hf00;
15'b0000101000101110111 : color = 12'hf11;
15'b0000101000101111000 : color = 12'hf73;
15'b0000101000101111001 : color = 12'he73;
15'b0000101000101111010 : color = 12'he73;
15'b0000101000101111011 : color = 12'he73;
15'b0000101000101111100 : color = 12'he73;
15'b0000101000101111101 : color = 12'he73;
15'b0000101000101111110 : color = 12'he73;
15'b0000101000101111111 : color = 12'he73;
15'b0000101000110000000 : color = 12'he73;
15'b0000101000110000001 : color = 12'he73;
15'b0000101000110000010 : color = 12'he73;
15'b0000101000110000011 : color = 12'he72;
15'b0000101000110000100 : color = 12'hf10;
15'b0000101000110000101 : color = 12'hf00;
15'b0000101000110000110 : color = 12'hf11;
15'b0000101000110000111 : color = 12'hf73;
15'b0000101000110001000 : color = 12'he73;
15'b0000101000110001001 : color = 12'he73;
15'b0000101000110001010 : color = 12'he73;
15'b0000101000110001011 : color = 12'he73;
15'b0000101000110001100 : color = 12'he73;
15'b0000101000110001101 : color = 12'he73;
15'b0000101000110001110 : color = 12'he73;
15'b0000101000110001111 : color = 12'he73;
15'b0000101000110010000 : color = 12'he73;
15'b0000101000110010001 : color = 12'he73;
15'b0000101000110010010 : color = 12'he73;
15'b0000101000110010011 : color = 12'he73;
15'b0000101000110010100 : color = 12'he73;
15'b0000101000110010101 : color = 12'he73;
15'b0000101000110010110 : color = 12'he73;
15'b0000101000110010111 : color = 12'he73;
15'b0000101000110011000 : color = 12'he73;
15'b0000101000110011001 : color = 12'he73;
15'b0000101000110011010 : color = 12'he73;
15'b0000101000110011011 : color = 12'he73;
15'b0000101000110011100 : color = 12'hf51;
15'b0000101000110011101 : color = 12'hf31;
15'b0000101000110011110 : color = 12'hf31;
15'b0000101000110011111 : color = 12'hf31;
15'b0000101000110100000 : color = 12'hf10;
15'b0000101000110100001 : color = 12'hf00;
15'b0000101000110100010 : color = 12'hf11;
15'b0000101000110100011 : color = 12'hf73;
15'b0000101000110100100 : color = 12'he73;
15'b0000101000110100101 : color = 12'hf30;
15'b0000101000110100110 : color = 12'hf11;
15'b0000101000110100111 : color = 12'hf73;
15'b0000101000110101000 : color = 12'he73;
15'b0000101000110101001 : color = 12'he73;
15'b0000101000110101010 : color = 12'he73;
15'b0000101000110101011 : color = 12'he61;
15'b0000101000110101100 : color = 12'hf00;
15'b0000101000110101101 : color = 12'hf53;
15'b0000101000110101110 : color = 12'he73;
15'b0000101000110101111 : color = 12'he73;
15'b0000101000110110000 : color = 12'he73;
15'b0000101000110110001 : color = 12'he73;
15'b0000101000110110010 : color = 12'he51;
15'b0000101000110110011 : color = 12'hf00;
15'b0000101000110110100 : color = 12'hf63;
15'b0000101000110110101 : color = 12'he73;
15'b0000101000110110110 : color = 12'he73;
15'b0000101000110110111 : color = 12'he73;
15'b0000101000110111000 : color = 12'he73;
15'b0000101000110111001 : color = 12'he73;
15'b0000101000110111010 : color = 12'he73;
15'b0000101000110111011 : color = 12'he73;
15'b0000101000110111100 : color = 12'he73;
15'b0000101000110111101 : color = 12'he73;
15'b0000101000110111110 : color = 12'he73;
15'b0000101000110111111 : color = 12'he73;
15'b0000101000111000000 : color = 12'he73;
15'b0000101000111000001 : color = 12'he73;
15'b0000101000111000010 : color = 12'he73;
15'b0000101000111000011 : color = 12'he73;
15'b0000101000111000100 : color = 12'he73;
15'b0000101000111000101 : color = 12'he73;
15'b0000101000111000110 : color = 12'he73;
15'b0000101000111000111 : color = 12'he73;
15'b0000101000111001000 : color = 12'he73;
15'b0000101000111001001 : color = 12'he51;
15'b0000101000111001010 : color = 12'hf01;
15'b0000101000111001011 : color = 12'hf73;
15'b0000101000111001100 : color = 12'he73;
15'b0000101000111001101 : color = 12'hf40;
15'b0000101000111001110 : color = 12'hf00;
15'b0000101000111001111 : color = 12'hf52;
15'b0000101000111010000 : color = 12'he73;
15'b0000101000111010001 : color = 12'he73;
15'b0000101000111010010 : color = 12'he73;
15'b0000101000111010011 : color = 12'he73;
15'b0000101000111010100 : color = 12'he73;
15'b0000101000111010101 : color = 12'he73;
15'b0000101000111010110 : color = 12'he73;
15'b0000101000111010111 : color = 12'he73;
15'b0000101000111011000 : color = 12'he73;
15'b0000101000111011001 : color = 12'he51;
15'b0000101000111011010 : color = 12'hf00;
15'b0000101000111011011 : color = 12'hf53;
15'b0000101000111011100 : color = 12'he73;
15'b0000101000111011101 : color = 12'he73;
15'b0000101000111011110 : color = 12'he73;
15'b0000101000111011111 : color = 12'he73;
15'b0000101000111100000 : color = 12'he73;
15'b0000101000111100001 : color = 12'he73;
15'b0000101000111100010 : color = 12'he73;
15'b0000101000111100011 : color = 12'he73;
15'b0000101000111100100 : color = 12'he73;
15'b0000101000111100101 : color = 12'he73;
15'b0000101000111100110 : color = 12'he73;
15'b0000101000111100111 : color = 12'he73;
15'b0000101000111101000 : color = 12'he73;
15'b0000101000111101001 : color = 12'he73;
15'b0000101000111101010 : color = 12'he73;
15'b0000101000111101011 : color = 12'he73;
15'b0000101000111101100 : color = 12'he73;
15'b0000101000111101101 : color = 12'he73;
15'b0000101000111101110 : color = 12'he73;
15'b0000101000111101111 : color = 12'he73;
15'b0000101000111110000 : color = 12'he73;
15'b0000101000111110001 : color = 12'he73;
15'b0000101000111110010 : color = 12'he73;
15'b0000101000111110011 : color = 12'he73;
15'b0000101000111110100 : color = 12'he73;
15'b0000101000111110101 : color = 12'he73;
15'b0000101000111110110 : color = 12'hf30;
15'b0000101000111110111 : color = 12'hf32;
15'b0000101000111111000 : color = 12'he73;
15'b0000101000111111001 : color = 12'he73;
15'b0000101000111111010 : color = 12'he73;
15'b0000101000111111011 : color = 12'he73;
15'b0000101000111111100 : color = 12'he73;
15'b0000101000111111101 : color = 12'he73;
15'b0000101000111111110 : color = 12'he73;
15'b0000101000111111111 : color = 12'he73;
15'b0000101001000000000 : color = 12'he73;
15'b0000101001000000001 : color = 12'he73;
15'b0000101001000000010 : color = 12'he73;
15'b0000101001000000011 : color = 12'he73;
15'b0000101001000000100 : color = 12'he73;
15'b0000101001000000101 : color = 12'he73;
15'b0000101001000000110 : color = 12'he73;
15'b0000101001000000111 : color = 12'he73;
15'b0000101001000001000 : color = 12'he73;
15'b0000101001000001001 : color = 12'he73;
15'b0000101001000001010 : color = 12'he72;
15'b0000101001000001011 : color = 12'hf10;
15'b0000101001000001100 : color = 12'hf00;
15'b0000101001000001101 : color = 12'hf42;
15'b0000101001000001110 : color = 12'hf73;
15'b0000101001000001111 : color = 12'he73;
15'b0000101001000010000 : color = 12'he73;
15'b0000101001000010001 : color = 12'he73;
15'b0000101001000010010 : color = 12'he73;
15'b0000101001000010011 : color = 12'he73;
15'b0000101001000010100 : color = 12'he73;
15'b0000101001000010101 : color = 12'he73;
15'b0000101001000010110 : color = 12'he73;
15'b0000101001000010111 : color = 12'he73;
15'b0000101001000011000 : color = 12'he73;
15'b0000101001000011001 : color = 12'he73;
15'b0000101001000011010 : color = 12'he73;
15'b0000101001000011011 : color = 12'he73;
15'b0000101001000011100 : color = 12'he73;
15'b0000101001000011101 : color = 12'he73;
15'b0000101001000011110 : color = 12'he73;
15'b0000101001000011111 : color = 12'he73;
15'b0000101001000100000 : color = 12'he73;
15'b0000101001000100001 : color = 12'he73;
15'b0000101001000100010 : color = 12'he73;
15'b0000101001000100011 : color = 12'he73;
15'b0000101001000100100 : color = 12'he72;
15'b0000101001000100101 : color = 12'hf10;
15'b0000101001000100110 : color = 12'hf32;
15'b0000101001000100111 : color = 12'he73;
15'b0000101001000101000 : color = 12'he73;
15'b0000101001000101001 : color = 12'he73;
15'b0000101001000101010 : color = 12'he73;
15'b0000101001000101011 : color = 12'he61;
15'b0000101001000101100 : color = 12'hf00;
15'b0000101001000101101 : color = 12'hf63;
15'b0000101001000101110 : color = 12'he73;
15'b0000101001000101111 : color = 12'he73;
15'b0000101001000110000 : color = 12'he73;
15'b0000101001000110001 : color = 12'hf30;
15'b0000101001000110010 : color = 12'hf32;
15'b0000101001000110011 : color = 12'he73;
15'b0000101001000110100 : color = 12'he73;
15'b0000101001000110101 : color = 12'he73;
15'b0000101001000110110 : color = 12'he61;
15'b0000101001000110111 : color = 12'hf00;
15'b0000101001000111000 : color = 12'hf63;
15'b0000101001000111001 : color = 12'he73;
15'b0000101001000111010 : color = 12'he73;
15'b0000101001000111011 : color = 12'he73;
15'b0000101001000111100 : color = 12'he73;
15'b0000101001000111101 : color = 12'he73;
15'b0000101001000111110 : color = 12'he73;
15'b0000101001000111111 : color = 12'he73;
15'b0000101001001000000 : color = 12'he73;
15'b0000101001001000001 : color = 12'he73;
15'b0000101001001000010 : color = 12'he73;
15'b0000101001001000011 : color = 12'he73;
15'b0000101001001000100 : color = 12'he73;
15'b0000101001001000101 : color = 12'he73;
15'b0000101001001000110 : color = 12'he73;
15'b0000101001001000111 : color = 12'he73;
15'b0000101001001001000 : color = 12'he73;
15'b0000101001001001001 : color = 12'he73;
15'b0000101001001001010 : color = 12'he73;
15'b0000101001001001011 : color = 12'he73;
15'b0000101001001001100 : color = 12'he73;
15'b0000101001001001101 : color = 12'he73;
15'b0000101001001001110 : color = 12'he73;
15'b0000101001001001111 : color = 12'he73;
15'b0000101001001010000 : color = 12'he73;
15'b0000101001001010001 : color = 12'he61;
15'b0000101001001010010 : color = 12'hf00;
15'b0000101001001010011 : color = 12'hf00;
15'b0000101001001010100 : color = 12'hf11;
15'b0000101001001010101 : color = 12'hf52;
15'b0000101001001010110 : color = 12'hf62;
15'b0000101001001010111 : color = 12'hf73;
15'b0000101001001011000 : color = 12'he73;
15'b0000101001001011001 : color = 12'he72;
15'b0000101001001011010 : color = 12'hf30;
15'b0000101001001011011 : color = 12'hf00;
15'b0000101001001011100 : color = 12'hf42;
15'b0000101001001011101 : color = 12'hf73;
15'b0000101001001011110 : color = 12'he73;
15'b0000101001001011111 : color = 12'he73;
15'b0000101001001100000 : color = 12'he73;
15'b0000101001001100001 : color = 12'he73;
15'b0000101001001100010 : color = 12'he73;
15'b0000101001001100011 : color = 12'he73;
15'b0000101001001100100 : color = 12'he73;
15'b0000101001001100101 : color = 12'he73;
15'b0000101001001100110 : color = 12'he73;
15'b0000101001001100111 : color = 12'he73;
15'b0000101001001101000 : color = 12'he73;
15'b0000101001001101001 : color = 12'he73;
15'b0000101001001101010 : color = 12'he73;
15'b0000101001001101011 : color = 12'he73;
15'b0000101001001101100 : color = 12'he73;
15'b0000101001001101101 : color = 12'he73;
15'b0000101001001101110 : color = 12'he73;
15'b0000101001001101111 : color = 12'he73;
15'b0000101001001110000 : color = 12'he73;
15'b0000101001001110001 : color = 12'he73;
15'b0000101001001110010 : color = 12'he73;
15'b0000101001001110011 : color = 12'he73;
15'b0000101001001110100 : color = 12'he73;
15'b0000101001001110101 : color = 12'he73;
15'b0000101001001110110 : color = 12'he73;
15'b0000101001001110111 : color = 12'he73;
15'b0000101001001111000 : color = 12'he73;
15'b0000101001001111001 : color = 12'hf40;
15'b0000101001001111010 : color = 12'hf11;
15'b0000101001001111011 : color = 12'hf52;
15'b0000101001001111100 : color = 12'hf73;
15'b0000101001001111101 : color = 12'he73;
15'b0000101001001111110 : color = 12'hf40;
15'b0000101001001111111 : color = 12'hf00;
15'b0000101001010000000 : color = 12'hf63;
15'b0000101001010000001 : color = 12'he73;
15'b0000101001010000010 : color = 12'he73;
15'b0000101001010000011 : color = 12'he73;
15'b0000101001010000100 : color = 12'he72;
15'b0000101001010000101 : color = 12'hf10;
15'b0000101001010000110 : color = 12'hf63;
15'b0000101001010000111 : color = 12'he73;
15'b0000101001010001000 : color = 12'he73;
15'b0000101001010001001 : color = 12'he73;
15'b0000101001010001010 : color = 12'he73;
15'b0000101001010001011 : color = 12'he73;
15'b0000101001010001100 : color = 12'he73;
15'b0000101001010001101 : color = 12'hf51;
15'b0000101001010001110 : color = 12'hf00;
15'b0000101001010001111 : color = 12'hf11;
15'b0000101001010010000 : color = 12'hf63;
15'b0000101001010010001 : color = 12'he73;
15'b0000101001010010010 : color = 12'he73;
15'b0000101001010010011 : color = 12'he73;
15'b0000101001010010100 : color = 12'he73;
15'b0000101001010010101 : color = 12'he73;
15'b0000101001010010110 : color = 12'he73;
15'b0000101001010010111 : color = 12'he73;
15'b0000101001010011000 : color = 12'he73;
15'b0000101001010011001 : color = 12'he73;
15'b0000101001010011010 : color = 12'he73;
15'b0000101001010011011 : color = 12'he73;
15'b0000101001010011100 : color = 12'he73;
15'b0000101001010011101 : color = 12'he73;
15'b0000101001010011110 : color = 12'he73;
15'b0000101001010011111 : color = 12'he73;
15'b0000101001010100000 : color = 12'he73;
15'b0000101001010100001 : color = 12'he73;
15'b0000101001010100010 : color = 12'he73;
15'b0000101000011100001 : color = 12'he73;
15'b0000101000011100010 : color = 12'he73;
15'b0000101000011100011 : color = 12'he73;
15'b0000101000011100100 : color = 12'he73;
15'b0000101000011100101 : color = 12'he73;
15'b0000101000011100110 : color = 12'he73;
15'b0000101000011100111 : color = 12'he73;
15'b0000101000011101000 : color = 12'he73;
15'b0000101000011101001 : color = 12'he73;
15'b0000101000011101010 : color = 12'he73;
15'b0000101000011101011 : color = 12'he73;
15'b0000101000011101100 : color = 12'he73;
15'b0000101000011101101 : color = 12'hf40;
15'b0000101000011101110 : color = 12'hf11;
15'b0000101000011101111 : color = 12'hf72;
15'b0000101000011110000 : color = 12'hf10;
15'b0000101000011110001 : color = 12'hf11;
15'b0000101000011110010 : color = 12'hf73;
15'b0000101000011110011 : color = 12'he73;
15'b0000101000011110100 : color = 12'he73;
15'b0000101000011110101 : color = 12'he51;
15'b0000101000011110110 : color = 12'hf42;
15'b0000101000011110111 : color = 12'he73;
15'b0000101000011111000 : color = 12'he73;
15'b0000101000011111001 : color = 12'he72;
15'b0000101000011111010 : color = 12'hf00;
15'b0000101000011111011 : color = 12'hf00;
15'b0000101000011111100 : color = 12'hf63;
15'b0000101000011111101 : color = 12'he73;
15'b0000101000011111110 : color = 12'he72;
15'b0000101000011111111 : color = 12'hf52;
15'b0000101000100000000 : color = 12'he73;
15'b0000101000100000001 : color = 12'he73;
15'b0000101000100000010 : color = 12'he73;
15'b0000101000100000011 : color = 12'he73;
15'b0000101000100000100 : color = 12'he73;
15'b0000101000100000101 : color = 12'he73;
15'b0000101000100000110 : color = 12'he73;
15'b0000101000100000111 : color = 12'he73;
15'b0000101000100001000 : color = 12'he73;
15'b0000101000100001001 : color = 12'he73;
15'b0000101000100001010 : color = 12'he73;
15'b0000101000100001011 : color = 12'he73;
15'b0000101000100001100 : color = 12'he73;
15'b0000101000100001101 : color = 12'he73;
15'b0000101000100001110 : color = 12'he73;
15'b0000101000100001111 : color = 12'he73;
15'b0000101000100010000 : color = 12'he73;
15'b0000101000100010001 : color = 12'he73;
15'b0000101000100010010 : color = 12'he73;
15'b0000101000100010011 : color = 12'he73;
15'b0000101000100010100 : color = 12'he73;
15'b0000101000100010101 : color = 12'he73;
15'b0000101000100010110 : color = 12'hf62;
15'b0000101000100010111 : color = 12'hf73;
15'b0000101000100011000 : color = 12'he73;
15'b0000101000100011001 : color = 12'he51;
15'b0000101000100011010 : color = 12'hf00;
15'b0000101000100011011 : color = 12'hf63;
15'b0000101000100011100 : color = 12'he73;
15'b0000101000100011101 : color = 12'he73;
15'b0000101000100011110 : color = 12'he61;
15'b0000101000100011111 : color = 12'hf00;
15'b0000101000100100000 : color = 12'hf53;
15'b0000101000100100001 : color = 12'he73;
15'b0000101000100100010 : color = 12'he73;
15'b0000101000100100011 : color = 12'he73;
15'b0000101000100100100 : color = 12'he73;
15'b0000101000100100101 : color = 12'he72;
15'b0000101000100100110 : color = 12'hf10;
15'b0000101000100100111 : color = 12'hf32;
15'b0000101000100101000 : color = 12'he73;
15'b0000101000100101001 : color = 12'he73;
15'b0000101000100101010 : color = 12'he73;
15'b0000101000100101011 : color = 12'he72;
15'b0000101000100101100 : color = 12'hf10;
15'b0000101000100101101 : color = 12'hf32;
15'b0000101000100101110 : color = 12'he73;
15'b0000101000100101111 : color = 12'he73;
15'b0000101000100110000 : color = 12'he73;
15'b0000101000100110001 : color = 12'he73;
15'b0000101000100110010 : color = 12'he73;
15'b0000101000100110011 : color = 12'he73;
15'b0000101000100110100 : color = 12'he73;
15'b0000101000100110101 : color = 12'he73;
15'b0000101000100110110 : color = 12'he73;
15'b0000101000100110111 : color = 12'he73;
15'b0000101000100111000 : color = 12'he73;
15'b0000101000100111001 : color = 12'he73;
15'b0000101000100111010 : color = 12'he73;
15'b0000101000100111011 : color = 12'he73;
15'b0000101000100111100 : color = 12'he73;
15'b0000101000100111101 : color = 12'he73;
15'b0000101000100111110 : color = 12'he73;
15'b0000101000100111111 : color = 12'he73;
15'b0000101000101000000 : color = 12'he73;
15'b0000101000101000001 : color = 12'he73;
15'b0000101000101000010 : color = 12'he73;
15'b0000101000101000011 : color = 12'he73;
15'b0000101000101000100 : color = 12'he73;
15'b0000101000101000101 : color = 12'he73;
15'b0000101000101000110 : color = 12'he73;
15'b0000101000101000111 : color = 12'he73;
15'b0000101000101001000 : color = 12'he51;
15'b0000101000101001001 : color = 12'hf00;
15'b0000101000101001010 : color = 12'hf53;
15'b0000101000101001011 : color = 12'he73;
15'b0000101000101001100 : color = 12'he73;
15'b0000101000101001101 : color = 12'he51;
15'b0000101000101001110 : color = 12'hf00;
15'b0000101000101001111 : color = 12'hf53;
15'b0000101000101010000 : color = 12'he73;
15'b0000101000101010001 : color = 12'he73;
15'b0000101000101010010 : color = 12'he51;
15'b0000101000101010011 : color = 12'hf01;
15'b0000101000101010100 : color = 12'hf63;
15'b0000101000101010101 : color = 12'he73;
15'b0000101000101010110 : color = 12'he73;
15'b0000101000101010111 : color = 12'he73;
15'b0000101000101011000 : color = 12'he73;
15'b0000101000101011001 : color = 12'hf63;
15'b0000101000101011010 : color = 12'he73;
15'b0000101000101011011 : color = 12'he73;
15'b0000101000101011100 : color = 12'he73;
15'b0000101000101011101 : color = 12'he73;
15'b0000101000101011110 : color = 12'he73;
15'b0000101000101011111 : color = 12'he73;
15'b0000101000101100000 : color = 12'he73;
15'b0000101000101100001 : color = 12'he73;
15'b0000101000101100010 : color = 12'he73;
15'b0000101000101100011 : color = 12'he73;
15'b0000101000101100100 : color = 12'he73;
15'b0000101000101100101 : color = 12'he73;
15'b0000101000101100110 : color = 12'he73;
15'b0000101000101100111 : color = 12'he73;
15'b0000101000101101000 : color = 12'he73;
15'b0000101000101101001 : color = 12'he73;
15'b0000101000101101010 : color = 12'he73;
15'b0000101000101101011 : color = 12'he73;
15'b0000101000101101100 : color = 12'he73;
15'b0000101000101101101 : color = 12'he73;
15'b0000101000101101110 : color = 12'he73;
15'b0000101000101101111 : color = 12'he51;
15'b0000101000101110000 : color = 12'hf00;
15'b0000101000101110001 : color = 12'hf10;
15'b0000101000101110010 : color = 12'hf31;
15'b0000101000101110011 : color = 12'hf52;
15'b0000101000101110100 : color = 12'hf62;
15'b0000101000101110101 : color = 12'hf00;
15'b0000101000101110110 : color = 12'hf42;
15'b0000101000101110111 : color = 12'he73;
15'b0000101000101111000 : color = 12'he73;
15'b0000101000101111001 : color = 12'he73;
15'b0000101000101111010 : color = 12'he61;
15'b0000101000101111011 : color = 12'hf00;
15'b0000101000101111100 : color = 12'hf01;
15'b0000101000101111101 : color = 12'hf73;
15'b0000101000101111110 : color = 12'he72;
15'b0000101000101111111 : color = 12'hf10;
15'b0000101000110000000 : color = 12'hf32;
15'b0000101000110000001 : color = 12'he73;
15'b0000101000110000010 : color = 12'he73;
15'b0000101000110000011 : color = 12'he73;
15'b0000101000110000100 : color = 12'hf40;
15'b0000101000110000101 : color = 12'hf01;
15'b0000101000110000110 : color = 12'hf73;
15'b0000101000110000111 : color = 12'he73;
15'b0000101000110001000 : color = 12'he73;
15'b0000101000110001001 : color = 12'he73;
15'b0000101000110001010 : color = 12'he73;
15'b0000101000110001011 : color = 12'he73;
15'b0000101000110001100 : color = 12'he73;
15'b0000101000110001101 : color = 12'he73;
15'b0000101000110001110 : color = 12'he73;
15'b0000101000110001111 : color = 12'he73;
15'b0000101000110010000 : color = 12'he73;
15'b0000101000110010001 : color = 12'he73;
15'b0000101000110010010 : color = 12'he73;
15'b0000101000110010011 : color = 12'he73;
15'b0000101000110010100 : color = 12'he73;
15'b0000101000110010101 : color = 12'he73;
15'b0000101000110010110 : color = 12'he73;
15'b0000101000110010111 : color = 12'he73;
15'b0000101000110011000 : color = 12'he73;
15'b0000101000110011001 : color = 12'he73;
15'b0000101000110011010 : color = 12'he73;
15'b0000101000110011011 : color = 12'he73;
15'b0000101000110011100 : color = 12'he73;
15'b0000101000110011101 : color = 12'he61;
15'b0000101000110011110 : color = 12'hf00;
15'b0000101000110011111 : color = 12'hf32;
15'b0000101000110100000 : color = 12'hf73;
15'b0000101000110100001 : color = 12'hf52;
15'b0000101000110100010 : color = 12'hf73;
15'b0000101000110100011 : color = 12'he73;
15'b0000101000110100100 : color = 12'he73;
15'b0000101000110100101 : color = 12'he73;
15'b0000101000110100110 : color = 12'he73;
15'b0000101000110100111 : color = 12'he73;
15'b0000101000110101000 : color = 12'he73;
15'b0000101000110101001 : color = 12'he61;
15'b0000101000110101010 : color = 12'hf11;
15'b0000101000110101011 : color = 12'hf63;
15'b0000101000110101100 : color = 12'he73;
15'b0000101000110101101 : color = 12'he72;
15'b0000101000110101110 : color = 12'hf10;
15'b0000101000110101111 : color = 12'hf00;
15'b0000101000110110000 : color = 12'hf11;
15'b0000101000110110001 : color = 12'hf73;
15'b0000101000110110010 : color = 12'he73;
15'b0000101000110110011 : color = 12'he73;
15'b0000101000110110100 : color = 12'he73;
15'b0000101000110110101 : color = 12'he73;
15'b0000101000110110110 : color = 12'he73;
15'b0000101000110110111 : color = 12'he73;
15'b0000101000110111000 : color = 12'he73;
15'b0000101000110111001 : color = 12'he73;
15'b0000101000110111010 : color = 12'he73;
15'b0000101000110111011 : color = 12'he73;
15'b0000101000110111100 : color = 12'he73;
15'b0000101000110111101 : color = 12'he73;
15'b0000101000110111110 : color = 12'he73;
15'b0000101000110111111 : color = 12'he73;
15'b0000101000111000000 : color = 12'he73;
15'b0000101000111000001 : color = 12'he73;
15'b0000101000111000010 : color = 12'he73;
15'b0000101000111000011 : color = 12'he73;
15'b0000101000111000100 : color = 12'he73;
15'b0000101000111000101 : color = 12'he72;
15'b0000101000111000110 : color = 12'hf62;
15'b0000101000111000111 : color = 12'he73;
15'b0000101000111001000 : color = 12'he73;
15'b0000101000111001001 : color = 12'he51;
15'b0000101000111001010 : color = 12'hf00;
15'b0000101000111001011 : color = 12'hf63;
15'b0000101000111001100 : color = 12'he73;
15'b0000101000111001101 : color = 12'he73;
15'b0000101000111001110 : color = 12'hf30;
15'b0000101000111001111 : color = 12'hf00;
15'b0000101000111010000 : color = 12'hf31;
15'b0000101000111010001 : color = 12'hf31;
15'b0000101000111010010 : color = 12'hf31;
15'b0000101000111010011 : color = 12'hf31;
15'b0000101000111010100 : color = 12'hf30;
15'b0000101000111010101 : color = 12'hf00;
15'b0000101000111010110 : color = 12'hf11;
15'b0000101000111010111 : color = 12'hf31;
15'b0000101000111011000 : color = 12'hf31;
15'b0000101000111011001 : color = 12'hf31;
15'b0000101000111011010 : color = 12'hf31;
15'b0000101000111011011 : color = 12'hf10;
15'b0000101000111011100 : color = 12'hf00;
15'b0000101000111011101 : color = 12'hf63;
15'b0000101000111011110 : color = 12'he73;
15'b0000101000111011111 : color = 12'he73;
15'b0000101000111100000 : color = 12'he73;
15'b0000101000111100001 : color = 12'he73;
15'b0000101000111100010 : color = 12'he73;
15'b0000101000111100011 : color = 12'he73;
15'b0000101000111100100 : color = 12'he73;
15'b0000101000111100101 : color = 12'he73;
15'b0000101000111100110 : color = 12'he73;
15'b0000101000111100111 : color = 12'he73;
15'b0000101000111101000 : color = 12'he73;
15'b0000101000111101001 : color = 12'he73;
15'b0000101000111101010 : color = 12'he73;
15'b0000101000111101011 : color = 12'he73;
15'b0000101000111101100 : color = 12'he73;
15'b0000101000111101101 : color = 12'he73;
15'b0000101000111101110 : color = 12'he73;
15'b0000101000111101111 : color = 12'he73;
15'b0000101000111110000 : color = 12'he73;
15'b0000101000111110001 : color = 12'he72;
15'b0000101000111110010 : color = 12'hf00;
15'b0000101000111110011 : color = 12'hf11;
15'b0000101000111110100 : color = 12'hf73;
15'b0000101000111110101 : color = 12'he73;
15'b0000101000111110110 : color = 12'hf40;
15'b0000101000111110111 : color = 12'hf01;
15'b0000101000111111000 : color = 12'hf73;
15'b0000101000111111001 : color = 12'he73;
15'b0000101000111111010 : color = 12'he73;
15'b0000101000111111011 : color = 12'he73;
15'b0000101000111111100 : color = 12'he73;
15'b0000101000111111101 : color = 12'he73;
15'b0000101000111111110 : color = 12'he73;
15'b0000101000111111111 : color = 12'he73;
15'b0000101001000000000 : color = 12'he73;
15'b0000101001000000001 : color = 12'he73;
15'b0000101001000000010 : color = 12'he51;
15'b0000101001000000011 : color = 12'hf00;
15'b0000101001000000100 : color = 12'hf53;
15'b0000101001000000101 : color = 12'he73;
15'b0000101001000000110 : color = 12'he73;
15'b0000101001000000111 : color = 12'he73;
15'b0000101001000001000 : color = 12'he73;
15'b0000101001000001001 : color = 12'he73;
15'b0000101001000001010 : color = 12'he73;
15'b0000101001000001011 : color = 12'he73;
15'b0000101001000001100 : color = 12'he73;
15'b0000101001000001101 : color = 12'he73;
15'b0000101001000001110 : color = 12'he73;
15'b0000101001000001111 : color = 12'he73;
15'b0000101001000010000 : color = 12'he73;
15'b0000101001000010001 : color = 12'he73;
15'b0000101001000010010 : color = 12'he73;
15'b0000101001000010011 : color = 12'he73;
15'b0000101001000010100 : color = 12'he73;
15'b0000101001000010101 : color = 12'he73;
15'b0000101001000010110 : color = 12'he73;
15'b0000101001000010111 : color = 12'he73;
15'b0000101001000011000 : color = 12'he73;
15'b0000101001000011001 : color = 12'he73;
15'b0000101001000011010 : color = 12'he73;
15'b0000101001000011011 : color = 12'he73;
15'b0000101001000011100 : color = 12'he73;
15'b0000101001000011101 : color = 12'he73;
15'b0000101001000011110 : color = 12'hf40;
15'b0000101001000011111 : color = 12'hf00;
15'b0000101001000100000 : color = 12'hf42;
15'b0000101001000100001 : color = 12'he73;
15'b0000101001000100010 : color = 12'he73;
15'b0000101001000100011 : color = 12'hf62;
15'b0000101001000100100 : color = 12'hf73;
15'b0000101001000100101 : color = 12'he73;
15'b0000101001000100110 : color = 12'he73;
15'b0000101001000100111 : color = 12'he73;
15'b0000101001000101000 : color = 12'he73;
15'b0000101001000101001 : color = 12'he73;
15'b0000101001000101010 : color = 12'he73;
15'b0000101001000101011 : color = 12'he73;
15'b0000101001000101100 : color = 12'he73;
15'b0000101001000101101 : color = 12'he73;
15'b0000101001000101110 : color = 12'he73;
15'b0000101001000101111 : color = 12'he51;
15'b0000101001000110000 : color = 12'hf52;
15'b0000101001000110001 : color = 12'he73;
15'b0000101001000110010 : color = 12'he73;
15'b0000101001000110011 : color = 12'he61;
15'b0000101001000110100 : color = 12'hf11;
15'b0000101001000110101 : color = 12'hf73;
15'b0000101001000110110 : color = 12'he73;
15'b0000101001000110111 : color = 12'he73;
15'b0000101001000111000 : color = 12'he73;
15'b0000101001000111001 : color = 12'he73;
15'b0000101001000111010 : color = 12'he73;
15'b0000101001000111011 : color = 12'he73;
15'b0000101001000111100 : color = 12'he73;
15'b0000101001000111101 : color = 12'he73;
15'b0000101001000111110 : color = 12'he73;
15'b0000101001000111111 : color = 12'he73;
15'b0000101001001000000 : color = 12'he73;
15'b0000101001001000001 : color = 12'he73;
15'b0000101001001000010 : color = 12'he73;
15'b0000101001001000011 : color = 12'he73;
15'b0000101001001000100 : color = 12'he73;
15'b0000101001001000101 : color = 12'he73;
15'b0000101001001000110 : color = 12'he73;
15'b0000101001001000111 : color = 12'he73;
15'b0000101001001001000 : color = 12'he73;
15'b0000101001001001001 : color = 12'he73;
15'b0000101001001001010 : color = 12'he73;
15'b0000101001001001011 : color = 12'he73;
15'b0000101001001001100 : color = 12'he73;
15'b0000101001001001101 : color = 12'he72;
15'b0000101001001001110 : color = 12'hf10;
15'b0000101001001001111 : color = 12'hf32;
15'b0000101001001010000 : color = 12'he73;
15'b0000101001001010001 : color = 12'hf40;
15'b0000101001001010010 : color = 12'hf32;
15'b0000101001001010011 : color = 12'he73;
15'b0000101001001010100 : color = 12'he61;
15'b0000101001001010101 : color = 12'hf00;
15'b0000101001001010110 : color = 12'hf63;
15'b0000101001001010111 : color = 12'he73;
15'b0000101001001011000 : color = 12'he73;
15'b0000101001001011001 : color = 12'he73;
15'b0000101001001011010 : color = 12'hf30;
15'b0000101001001011011 : color = 12'hf32;
15'b0000101001001011100 : color = 12'he73;
15'b0000101001001011101 : color = 12'he73;
15'b0000101001001011110 : color = 12'he73;
15'b0000101001001011111 : color = 12'he61;
15'b0000101001001100000 : color = 12'hf00;
15'b0000101001001100001 : color = 12'hf63;
15'b0000101001001100010 : color = 12'he73;
15'b0000101001001100011 : color = 12'he73;
15'b0000101001001100100 : color = 12'he73;
15'b0000101001001100101 : color = 12'he73;
15'b0000101001001100110 : color = 12'he73;
15'b0000101001001100111 : color = 12'he73;
15'b0000101001001101000 : color = 12'he73;
15'b0000101001001101001 : color = 12'he73;
15'b0000101001001101010 : color = 12'he73;
15'b0000101001001101011 : color = 12'he73;
15'b0000101001001101100 : color = 12'he73;
15'b0000101001001101101 : color = 12'he73;
15'b0000101001001101110 : color = 12'he73;
15'b0000101001001101111 : color = 12'he73;
15'b0000101001001110000 : color = 12'he73;
15'b0000101001001110001 : color = 12'he73;
15'b0000101001001110010 : color = 12'he73;
15'b0000101001001110011 : color = 12'he73;
15'b0000101001001110100 : color = 12'he73;
15'b0000101001001110101 : color = 12'he73;
15'b0000101001001110110 : color = 12'he73;
15'b0000101001001110111 : color = 12'he73;
15'b0000101001001111000 : color = 12'he73;
15'b0000101001001111001 : color = 12'he73;
15'b0000101001001111010 : color = 12'he73;
15'b0000101001001111011 : color = 12'hf62;
15'b0000101001001111100 : color = 12'he73;
15'b0000101001001111101 : color = 12'he73;
15'b0000101001001111110 : color = 12'he73;
15'b0000101001001111111 : color = 12'he73;
15'b0000101001010000000 : color = 12'he73;
15'b0000101001010000001 : color = 12'hf51;
15'b0000101001010000010 : color = 12'hf00;
15'b0000101001010000011 : color = 12'hf32;
15'b0000101001010000100 : color = 12'hf73;
15'b0000101001010000101 : color = 12'he73;
15'b0000101001010000110 : color = 12'he73;
15'b0000101001010000111 : color = 12'he73;
15'b0000101001010001000 : color = 12'he73;
15'b0000101001010001001 : color = 12'he73;
15'b0000101001010001010 : color = 12'he73;
15'b0000101001010001011 : color = 12'he73;
15'b0000101001010001100 : color = 12'he73;
15'b0000101001010001101 : color = 12'he73;
15'b0000101001010001110 : color = 12'he73;
15'b0000101001010001111 : color = 12'he73;
15'b0000101001010010000 : color = 12'he73;
15'b0000101001010010001 : color = 12'he73;
15'b0000101001010010010 : color = 12'he73;
15'b0000101001010010011 : color = 12'he73;
15'b0000101001010010100 : color = 12'he73;
15'b0000101001010010101 : color = 12'he73;
15'b0000101001010010110 : color = 12'he73;
15'b0000101001010010111 : color = 12'he73;
15'b0000101001010011000 : color = 12'he73;
15'b0000101001010011001 : color = 12'he73;
15'b0000101001010011010 : color = 12'he73;
15'b0000101001010011011 : color = 12'he73;
15'b0000101001010011100 : color = 12'he73;
15'b0000101001010011101 : color = 12'he73;
15'b0000101001010011110 : color = 12'he73;
15'b0000101001010011111 : color = 12'he73;
15'b0000101001010100000 : color = 12'he73;
15'b0000101001010100001 : color = 12'he73;
15'b0000101001010100010 : color = 12'he73;
15'b0000101001010100011 : color = 12'he73;
15'b0000101001010100100 : color = 12'he73;
15'b0000101001010100101 : color = 12'he73;
15'b0000101001010100110 : color = 12'he61;
15'b0000101001010100111 : color = 12'hf00;
15'b0000101001010101000 : color = 12'hf53;
15'b0000101001010101001 : color = 12'he73;
15'b0000101001010101010 : color = 12'he73;
15'b0000101001010101011 : color = 12'he73;
15'b0000101001010101100 : color = 12'he62;
15'b0000101001010101101 : color = 12'hf10;
15'b0000101001010101110 : color = 12'hf52;
15'b0000101001010101111 : color = 12'hf62;
15'b0000101001010110000 : color = 12'hf62;
15'b0000101001010110001 : color = 12'hf62;
15'b0000101001010110010 : color = 12'hf62;
15'b0000101001010110011 : color = 12'hf52;
15'b0000101001010110100 : color = 12'hf52;
15'b0000101001010110101 : color = 12'hf52;
15'b0000101001010110110 : color = 12'hf51;
15'b0000101001010110111 : color = 12'hf10;
15'b0000101001010111000 : color = 12'hf00;
15'b0000101001010111001 : color = 12'hf01;
15'b0000101001010111010 : color = 12'hf73;
15'b0000101001010111011 : color = 12'he73;
15'b0000101001010111100 : color = 12'he73;
15'b0000101001010111101 : color = 12'he73;
15'b0000101001010111110 : color = 12'he73;
15'b0000101001010111111 : color = 12'he73;
15'b0000101001011000000 : color = 12'he73;
15'b0000101001011000001 : color = 12'he73;
15'b0000101001011000010 : color = 12'he73;
15'b0000101001011000011 : color = 12'he73;
15'b0000101001011000100 : color = 12'he73;
15'b0000101001011000101 : color = 12'he73;
15'b0000101001011000110 : color = 12'he73;
15'b0000101001011000111 : color = 12'he73;
15'b0000101001011001000 : color = 12'he73;
15'b0000101001011001001 : color = 12'he73;
15'b0000101001011001010 : color = 12'he73;
15'b0000101001011001011 : color = 12'he73;
15'b0000101000100001010 : color = 12'he73;
15'b0000101000100001011 : color = 12'he73;
15'b0000101000100001100 : color = 12'he73;
15'b0000101000100001101 : color = 12'he73;
15'b0000101000100001110 : color = 12'he73;
15'b0000101000100001111 : color = 12'he73;
15'b0000101000100010000 : color = 12'he73;
15'b0000101000100010001 : color = 12'he73;
15'b0000101000100010010 : color = 12'he73;
15'b0000101000100010011 : color = 12'he73;
15'b0000101000100010100 : color = 12'he73;
15'b0000101000100010101 : color = 12'he73;
15'b0000101000100010110 : color = 12'he72;
15'b0000101000100010111 : color = 12'hf10;
15'b0000101000100011000 : color = 12'hf10;
15'b0000101000100011001 : color = 12'hf00;
15'b0000101000100011010 : color = 12'hf53;
15'b0000101000100011011 : color = 12'he73;
15'b0000101000100011100 : color = 12'he73;
15'b0000101000100011101 : color = 12'he72;
15'b0000101000100011110 : color = 12'hf11;
15'b0000101000100011111 : color = 12'hf73;
15'b0000101000100100000 : color = 12'he73;
15'b0000101000100100001 : color = 12'he73;
15'b0000101000100100010 : color = 12'he61;
15'b0000101000100100011 : color = 12'hf00;
15'b0000101000100100100 : color = 12'hf31;
15'b0000101000100100101 : color = 12'hf53;
15'b0000101000100100110 : color = 12'he73;
15'b0000101000100100111 : color = 12'he73;
15'b0000101000100101000 : color = 12'he73;
15'b0000101000100101001 : color = 12'he73;
15'b0000101000100101010 : color = 12'he73;
15'b0000101000100101011 : color = 12'he73;
15'b0000101000100101100 : color = 12'he73;
15'b0000101000100101101 : color = 12'he73;
15'b0000101000100101110 : color = 12'he73;
15'b0000101000100101111 : color = 12'he73;
15'b0000101000100110000 : color = 12'he73;
15'b0000101000100110001 : color = 12'he73;
15'b0000101000100110010 : color = 12'he73;
15'b0000101000100110011 : color = 12'he73;
15'b0000101000100110100 : color = 12'he73;
15'b0000101000100110101 : color = 12'he73;
15'b0000101000100110110 : color = 12'he73;
15'b0000101000100110111 : color = 12'he73;
15'b0000101000100111000 : color = 12'he73;
15'b0000101000100111001 : color = 12'he73;
15'b0000101000100111010 : color = 12'he73;
15'b0000101000100111011 : color = 12'he73;
15'b0000101000100111100 : color = 12'he73;
15'b0000101000100111101 : color = 12'he73;
15'b0000101000100111110 : color = 12'he73;
15'b0000101000100111111 : color = 12'he73;
15'b0000101000101000000 : color = 12'he73;
15'b0000101000101000001 : color = 12'he73;
15'b0000101000101000010 : color = 12'he51;
15'b0000101000101000011 : color = 12'hf00;
15'b0000101000101000100 : color = 12'hf63;
15'b0000101000101000101 : color = 12'he73;
15'b0000101000101000110 : color = 12'he73;
15'b0000101000101000111 : color = 12'he61;
15'b0000101000101001000 : color = 12'hf00;
15'b0000101000101001001 : color = 12'hf53;
15'b0000101000101001010 : color = 12'he73;
15'b0000101000101001011 : color = 12'he73;
15'b0000101000101001100 : color = 12'he73;
15'b0000101000101001101 : color = 12'he73;
15'b0000101000101001110 : color = 12'he72;
15'b0000101000101001111 : color = 12'hf10;
15'b0000101000101010000 : color = 12'hf32;
15'b0000101000101010001 : color = 12'he73;
15'b0000101000101010010 : color = 12'he73;
15'b0000101000101010011 : color = 12'he73;
15'b0000101000101010100 : color = 12'he72;
15'b0000101000101010101 : color = 12'hf10;
15'b0000101000101010110 : color = 12'hf32;
15'b0000101000101010111 : color = 12'he73;
15'b0000101000101011000 : color = 12'he73;
15'b0000101000101011001 : color = 12'he73;
15'b0000101000101011010 : color = 12'he73;
15'b0000101000101011011 : color = 12'he73;
15'b0000101000101011100 : color = 12'he73;
15'b0000101000101011101 : color = 12'he73;
15'b0000101000101011110 : color = 12'he73;
15'b0000101000101011111 : color = 12'he73;
15'b0000101000101100000 : color = 12'he73;
15'b0000101000101100001 : color = 12'he73;
15'b0000101000101100010 : color = 12'he73;
15'b0000101000101100011 : color = 12'he73;
15'b0000101000101100100 : color = 12'he73;
15'b0000101000101100101 : color = 12'he73;
15'b0000101000101100110 : color = 12'he73;
15'b0000101000101100111 : color = 12'he73;
15'b0000101000101101000 : color = 12'he73;
15'b0000101000101101001 : color = 12'he73;
15'b0000101000101101010 : color = 12'he73;
15'b0000101000101101011 : color = 12'he73;
15'b0000101000101101100 : color = 12'he73;
15'b0000101000101101101 : color = 12'he73;
15'b0000101000101101110 : color = 12'he73;
15'b0000101000101101111 : color = 12'he73;
15'b0000101000101110000 : color = 12'he73;
15'b0000101000101110001 : color = 12'he72;
15'b0000101000101110010 : color = 12'hf31;
15'b0000101000101110011 : color = 12'hf73;
15'b0000101000101110100 : color = 12'he73;
15'b0000101000101110101 : color = 12'he73;
15'b0000101000101110110 : color = 12'he51;
15'b0000101000101110111 : color = 12'hf00;
15'b0000101000101111000 : color = 12'hf53;
15'b0000101000101111001 : color = 12'he73;
15'b0000101000101111010 : color = 12'he72;
15'b0000101000101111011 : color = 12'hf11;
15'b0000101000101111100 : color = 12'hf63;
15'b0000101000101111101 : color = 12'he73;
15'b0000101000101111110 : color = 12'he73;
15'b0000101000101111111 : color = 12'he73;
15'b0000101000110000000 : color = 12'he73;
15'b0000101000110000001 : color = 12'hf30;
15'b0000101000110000010 : color = 12'hf00;
15'b0000101000110000011 : color = 12'hf63;
15'b0000101000110000100 : color = 12'he73;
15'b0000101000110000101 : color = 12'he73;
15'b0000101000110000110 : color = 12'he73;
15'b0000101000110000111 : color = 12'he73;
15'b0000101000110001000 : color = 12'he73;
15'b0000101000110001001 : color = 12'he73;
15'b0000101000110001010 : color = 12'he73;
15'b0000101000110001011 : color = 12'he73;
15'b0000101000110001100 : color = 12'he73;
15'b0000101000110001101 : color = 12'he73;
15'b0000101000110001110 : color = 12'he73;
15'b0000101000110001111 : color = 12'he73;
15'b0000101000110010000 : color = 12'he73;
15'b0000101000110010001 : color = 12'he73;
15'b0000101000110010010 : color = 12'he73;
15'b0000101000110010011 : color = 12'he73;
15'b0000101000110010100 : color = 12'he73;
15'b0000101000110010101 : color = 12'he73;
15'b0000101000110010110 : color = 12'he73;
15'b0000101000110010111 : color = 12'he73;
15'b0000101000110011000 : color = 12'he73;
15'b0000101000110011001 : color = 12'hf63;
15'b0000101000110011010 : color = 12'he73;
15'b0000101000110011011 : color = 12'he73;
15'b0000101000110011100 : color = 12'he73;
15'b0000101000110011101 : color = 12'he72;
15'b0000101000110011110 : color = 12'hf00;
15'b0000101000110011111 : color = 12'hf11;
15'b0000101000110100000 : color = 12'hf73;
15'b0000101000110100001 : color = 12'he73;
15'b0000101000110100010 : color = 12'he73;
15'b0000101000110100011 : color = 12'he73;
15'b0000101000110100100 : color = 12'hf30;
15'b0000101000110100101 : color = 12'hf32;
15'b0000101000110100110 : color = 12'hf73;
15'b0000101000110100111 : color = 12'he72;
15'b0000101000110101000 : color = 12'hf10;
15'b0000101000110101001 : color = 12'hf32;
15'b0000101000110101010 : color = 12'he73;
15'b0000101000110101011 : color = 12'he73;
15'b0000101000110101100 : color = 12'he73;
15'b0000101000110101101 : color = 12'hf40;
15'b0000101000110101110 : color = 12'hf01;
15'b0000101000110101111 : color = 12'hf73;
15'b0000101000110110000 : color = 12'he73;
15'b0000101000110110001 : color = 12'he73;
15'b0000101000110110010 : color = 12'he73;
15'b0000101000110110011 : color = 12'he73;
15'b0000101000110110100 : color = 12'he73;
15'b0000101000110110101 : color = 12'he73;
15'b0000101000110110110 : color = 12'he73;
15'b0000101000110110111 : color = 12'he73;
15'b0000101000110111000 : color = 12'he73;
15'b0000101000110111001 : color = 12'he73;
15'b0000101000110111010 : color = 12'he73;
15'b0000101000110111011 : color = 12'he73;
15'b0000101000110111100 : color = 12'he73;
15'b0000101000110111101 : color = 12'he73;
15'b0000101000110111110 : color = 12'he73;
15'b0000101000110111111 : color = 12'he73;
15'b0000101000111000000 : color = 12'he73;
15'b0000101000111000001 : color = 12'he73;
15'b0000101000111000010 : color = 12'he73;
15'b0000101000111000011 : color = 12'he73;
15'b0000101000111000100 : color = 12'he73;
15'b0000101000111000101 : color = 12'hf51;
15'b0000101000111000110 : color = 12'hf00;
15'b0000101000111000111 : color = 12'hf52;
15'b0000101000111001000 : color = 12'he73;
15'b0000101000111001001 : color = 12'he73;
15'b0000101000111001010 : color = 12'he51;
15'b0000101000111001011 : color = 12'hf63;
15'b0000101000111001100 : color = 12'he73;
15'b0000101000111001101 : color = 12'he73;
15'b0000101000111001110 : color = 12'he73;
15'b0000101000111001111 : color = 12'he73;
15'b0000101000111010000 : color = 12'he73;
15'b0000101000111010001 : color = 12'he73;
15'b0000101000111010010 : color = 12'hf40;
15'b0000101000111010011 : color = 12'hf00;
15'b0000101000111010100 : color = 12'hf00;
15'b0000101000111010101 : color = 12'hf52;
15'b0000101000111010110 : color = 12'he73;
15'b0000101000111010111 : color = 12'he72;
15'b0000101000111011000 : color = 12'hf00;
15'b0000101000111011001 : color = 12'hf01;
15'b0000101000111011010 : color = 12'hf73;
15'b0000101000111011011 : color = 12'he73;
15'b0000101000111011100 : color = 12'he73;
15'b0000101000111011101 : color = 12'he73;
15'b0000101000111011110 : color = 12'he73;
15'b0000101000111011111 : color = 12'he73;
15'b0000101000111100000 : color = 12'he73;
15'b0000101000111100001 : color = 12'he73;
15'b0000101000111100010 : color = 12'he73;
15'b0000101000111100011 : color = 12'he73;
15'b0000101000111100100 : color = 12'he73;
15'b0000101000111100101 : color = 12'he73;
15'b0000101000111100110 : color = 12'he73;
15'b0000101000111100111 : color = 12'he73;
15'b0000101000111101000 : color = 12'he73;
15'b0000101000111101001 : color = 12'he73;
15'b0000101000111101010 : color = 12'he73;
15'b0000101000111101011 : color = 12'he73;
15'b0000101000111101100 : color = 12'he73;
15'b0000101000111101101 : color = 12'he73;
15'b0000101000111101110 : color = 12'he73;
15'b0000101000111101111 : color = 12'he73;
15'b0000101000111110000 : color = 12'he73;
15'b0000101000111110001 : color = 12'he73;
15'b0000101000111110010 : color = 12'he51;
15'b0000101000111110011 : color = 12'hf00;
15'b0000101000111110100 : color = 12'hf63;
15'b0000101000111110101 : color = 12'he73;
15'b0000101000111110110 : color = 12'he73;
15'b0000101000111110111 : color = 12'hf40;
15'b0000101000111111000 : color = 12'hf11;
15'b0000101000111111001 : color = 12'hf73;
15'b0000101000111111010 : color = 12'he73;
15'b0000101000111111011 : color = 12'he73;
15'b0000101000111111100 : color = 12'he73;
15'b0000101000111111101 : color = 12'he61;
15'b0000101000111111110 : color = 12'hf00;
15'b0000101000111111111 : color = 12'hf53;
15'b0000101001000000000 : color = 12'he73;
15'b0000101001000000001 : color = 12'he73;
15'b0000101001000000010 : color = 12'he73;
15'b0000101001000000011 : color = 12'he73;
15'b0000101001000000100 : color = 12'he51;
15'b0000101001000000101 : color = 12'hf00;
15'b0000101001000000110 : color = 12'hf63;
15'b0000101001000000111 : color = 12'he73;
15'b0000101001000001000 : color = 12'he73;
15'b0000101001000001001 : color = 12'he73;
15'b0000101001000001010 : color = 12'he73;
15'b0000101001000001011 : color = 12'he73;
15'b0000101001000001100 : color = 12'he73;
15'b0000101001000001101 : color = 12'he73;
15'b0000101001000001110 : color = 12'he73;
15'b0000101001000001111 : color = 12'he73;
15'b0000101001000010000 : color = 12'he73;
15'b0000101001000010001 : color = 12'he73;
15'b0000101001000010010 : color = 12'he73;
15'b0000101001000010011 : color = 12'he73;
15'b0000101001000010100 : color = 12'he73;
15'b0000101001000010101 : color = 12'he73;
15'b0000101001000010110 : color = 12'he73;
15'b0000101001000010111 : color = 12'he73;
15'b0000101001000011000 : color = 12'he73;
15'b0000101001000011001 : color = 12'he73;
15'b0000101001000011010 : color = 12'hf30;
15'b0000101001000011011 : color = 12'hf00;
15'b0000101001000011100 : color = 12'hf42;
15'b0000101001000011101 : color = 12'he73;
15'b0000101001000011110 : color = 12'he73;
15'b0000101001000011111 : color = 12'hf40;
15'b0000101001000100000 : color = 12'hf01;
15'b0000101001000100001 : color = 12'hf73;
15'b0000101001000100010 : color = 12'he73;
15'b0000101001000100011 : color = 12'he73;
15'b0000101001000100100 : color = 12'he73;
15'b0000101001000100101 : color = 12'he73;
15'b0000101001000100110 : color = 12'he73;
15'b0000101001000100111 : color = 12'he73;
15'b0000101001000101000 : color = 12'he73;
15'b0000101001000101001 : color = 12'he73;
15'b0000101001000101010 : color = 12'he73;
15'b0000101001000101011 : color = 12'he51;
15'b0000101001000101100 : color = 12'hf00;
15'b0000101001000101101 : color = 12'hf53;
15'b0000101001000101110 : color = 12'he73;
15'b0000101001000101111 : color = 12'he73;
15'b0000101001000110000 : color = 12'he73;
15'b0000101001000110001 : color = 12'he73;
15'b0000101001000110010 : color = 12'he73;
15'b0000101001000110011 : color = 12'he73;
15'b0000101001000110100 : color = 12'he73;
15'b0000101001000110101 : color = 12'he73;
15'b0000101001000110110 : color = 12'he73;
15'b0000101001000110111 : color = 12'he73;
15'b0000101001000111000 : color = 12'he73;
15'b0000101001000111001 : color = 12'he73;
15'b0000101001000111010 : color = 12'he73;
15'b0000101001000111011 : color = 12'he73;
15'b0000101001000111100 : color = 12'he73;
15'b0000101001000111101 : color = 12'he73;
15'b0000101001000111110 : color = 12'he73;
15'b0000101001000111111 : color = 12'he73;
15'b0000101001001000000 : color = 12'he73;
15'b0000101001001000001 : color = 12'he73;
15'b0000101001001000010 : color = 12'he73;
15'b0000101001001000011 : color = 12'he73;
15'b0000101001001000100 : color = 12'he73;
15'b0000101001001000101 : color = 12'he73;
15'b0000101001001000110 : color = 12'he62;
15'b0000101001001000111 : color = 12'hf00;
15'b0000101001001001000 : color = 12'hf11;
15'b0000101001001001001 : color = 12'hf73;
15'b0000101001001001010 : color = 12'he73;
15'b0000101001001001011 : color = 12'he73;
15'b0000101001001001100 : color = 12'hf30;
15'b0000101001001001101 : color = 12'hf10;
15'b0000101001001001110 : color = 12'hf31;
15'b0000101001001001111 : color = 12'hf31;
15'b0000101001001010000 : color = 12'hf31;
15'b0000101001001010001 : color = 12'hf31;
15'b0000101001001010010 : color = 12'hf31;
15'b0000101001001010011 : color = 12'hf31;
15'b0000101001001010100 : color = 12'hf31;
15'b0000101001001010101 : color = 12'hf31;
15'b0000101001001010110 : color = 12'hf31;
15'b0000101001001010111 : color = 12'hf31;
15'b0000101001001011000 : color = 12'hf00;
15'b0000101001001011001 : color = 12'hf00;
15'b0000101001001011010 : color = 12'hf53;
15'b0000101001001011011 : color = 12'he73;
15'b0000101001001011100 : color = 12'hf41;
15'b0000101001001011101 : color = 12'hf73;
15'b0000101001001011110 : color = 12'he73;
15'b0000101001001011111 : color = 12'he73;
15'b0000101001001100000 : color = 12'he73;
15'b0000101001001100001 : color = 12'he73;
15'b0000101001001100010 : color = 12'he73;
15'b0000101001001100011 : color = 12'he73;
15'b0000101001001100100 : color = 12'he73;
15'b0000101001001100101 : color = 12'he73;
15'b0000101001001100110 : color = 12'he73;
15'b0000101001001100111 : color = 12'he73;
15'b0000101001001101000 : color = 12'he73;
15'b0000101001001101001 : color = 12'he73;
15'b0000101001001101010 : color = 12'he73;
15'b0000101001001101011 : color = 12'he73;
15'b0000101001001101100 : color = 12'he73;
15'b0000101001001101101 : color = 12'he73;
15'b0000101001001101110 : color = 12'he73;
15'b0000101001001101111 : color = 12'he73;
15'b0000101001001110000 : color = 12'he73;
15'b0000101001001110001 : color = 12'he73;
15'b0000101001001110010 : color = 12'he72;
15'b0000101001001110011 : color = 12'hf41;
15'b0000101001001110100 : color = 12'hf31;
15'b0000101001001110101 : color = 12'hf31;
15'b0000101001001110110 : color = 12'hf31;
15'b0000101001001110111 : color = 12'hf00;
15'b0000101001001111000 : color = 12'hf10;
15'b0000101001001111001 : color = 12'hf30;
15'b0000101001001111010 : color = 12'hf00;
15'b0000101001001111011 : color = 12'hf00;
15'b0000101001001111100 : color = 12'hf42;
15'b0000101001001111101 : color = 12'he61;
15'b0000101001001111110 : color = 12'hf00;
15'b0000101001001111111 : color = 12'hf63;
15'b0000101001010000000 : color = 12'he73;
15'b0000101001010000001 : color = 12'he73;
15'b0000101001010000010 : color = 12'he73;
15'b0000101001010000011 : color = 12'hf30;
15'b0000101001010000100 : color = 12'hf32;
15'b0000101001010000101 : color = 12'he73;
15'b0000101001010000110 : color = 12'he73;
15'b0000101001010000111 : color = 12'he73;
15'b0000101001010001000 : color = 12'he61;
15'b0000101001010001001 : color = 12'hf00;
15'b0000101001010001010 : color = 12'hf63;
15'b0000101001010001011 : color = 12'he73;
15'b0000101001010001100 : color = 12'he73;
15'b0000101001010001101 : color = 12'he73;
15'b0000101001010001110 : color = 12'he73;
15'b0000101001010001111 : color = 12'he73;
15'b0000101001010010000 : color = 12'he73;
15'b0000101001010010001 : color = 12'he73;
15'b0000101001010010010 : color = 12'he73;
15'b0000101001010010011 : color = 12'he73;
15'b0000101001010010100 : color = 12'he73;
15'b0000101001010010101 : color = 12'he73;
15'b0000101001010010110 : color = 12'he73;
15'b0000101001010010111 : color = 12'he73;
15'b0000101001010011000 : color = 12'he73;
15'b0000101001010011001 : color = 12'he73;
15'b0000101001010011010 : color = 12'he73;
15'b0000101001010011011 : color = 12'he73;
15'b0000101001010011100 : color = 12'he73;
15'b0000101001010011101 : color = 12'he73;
15'b0000101001010011110 : color = 12'he73;
15'b0000101001010011111 : color = 12'he73;
15'b0000101001010100000 : color = 12'he73;
15'b0000101001010100001 : color = 12'he73;
15'b0000101001010100010 : color = 12'he73;
15'b0000101001010100011 : color = 12'he73;
15'b0000101001010100100 : color = 12'he73;
15'b0000101001010100101 : color = 12'he73;
15'b0000101001010100110 : color = 12'he73;
15'b0000101001010100111 : color = 12'he73;
15'b0000101001010101000 : color = 12'hf51;
15'b0000101001010101001 : color = 12'hf10;
15'b0000101001010101010 : color = 12'hf11;
15'b0000101001010101011 : color = 12'hf63;
15'b0000101001010101100 : color = 12'he73;
15'b0000101001010101101 : color = 12'he73;
15'b0000101001010101110 : color = 12'he73;
15'b0000101001010101111 : color = 12'he73;
15'b0000101001010110000 : color = 12'he51;
15'b0000101001010110001 : color = 12'hf11;
15'b0000101001010110010 : color = 12'hf52;
15'b0000101001010110011 : color = 12'he73;
15'b0000101001010110100 : color = 12'he73;
15'b0000101001010110101 : color = 12'he73;
15'b0000101001010110110 : color = 12'he73;
15'b0000101001010110111 : color = 12'he73;
15'b0000101001010111000 : color = 12'he73;
15'b0000101001010111001 : color = 12'he73;
15'b0000101001010111010 : color = 12'he73;
15'b0000101001010111011 : color = 12'he73;
15'b0000101001010111100 : color = 12'he73;
15'b0000101001010111101 : color = 12'he73;
15'b0000101001010111110 : color = 12'he73;
15'b0000101001010111111 : color = 12'he73;
15'b0000101001011000000 : color = 12'he73;
15'b0000101001011000001 : color = 12'he73;
15'b0000101001011000010 : color = 12'he73;
15'b0000101001011000011 : color = 12'he73;
15'b0000101001011000100 : color = 12'he73;
15'b0000101001011000101 : color = 12'he73;
15'b0000101001011000110 : color = 12'he73;
15'b0000101001011000111 : color = 12'he73;
15'b0000101001011001000 : color = 12'he73;
15'b0000101001011001001 : color = 12'he73;
15'b0000101001011001010 : color = 12'he73;
15'b0000101001011001011 : color = 12'he73;
15'b0000101001011001100 : color = 12'he73;
15'b0000101001011001101 : color = 12'he73;
15'b0000101001011001110 : color = 12'he72;
15'b0000101001011001111 : color = 12'hf00;
15'b0000101001011010000 : color = 12'hf42;
15'b0000101001011010001 : color = 12'he73;
15'b0000101001011010010 : color = 12'he73;
15'b0000101001011010011 : color = 12'he73;
15'b0000101001011010100 : color = 12'he73;
15'b0000101001011010101 : color = 12'hf30;
15'b0000101001011010110 : color = 12'hf00;
15'b0000101001011010111 : color = 12'hf00;
15'b0000101001011011000 : color = 12'hf00;
15'b0000101001011011001 : color = 12'hf00;
15'b0000101001011011010 : color = 12'hf10;
15'b0000101001011011011 : color = 12'hf31;
15'b0000101001011011100 : color = 12'hf41;
15'b0000101001011011101 : color = 12'hf51;
15'b0000101001011011110 : color = 12'hf52;
15'b0000101001011011111 : color = 12'hf62;
15'b0000101001011100000 : color = 12'he73;
15'b0000101001011100001 : color = 12'hf30;
15'b0000101001011100010 : color = 12'hf00;
15'b0000101001011100011 : color = 12'hf63;
15'b0000101001011100100 : color = 12'he73;
15'b0000101001011100101 : color = 12'he73;
15'b0000101001011100110 : color = 12'he73;
15'b0000101001011100111 : color = 12'he73;
15'b0000101001011101000 : color = 12'he73;
15'b0000101001011101001 : color = 12'he73;
15'b0000101001011101010 : color = 12'he73;
15'b0000101001011101011 : color = 12'he73;
15'b0000101001011101100 : color = 12'he73;
15'b0000101001011101101 : color = 12'he73;
15'b0000101001011101110 : color = 12'he73;
15'b0000101001011101111 : color = 12'he73;
15'b0000101001011110000 : color = 12'he73;
15'b0000101001011110001 : color = 12'he73;
15'b0000101001011110010 : color = 12'he73;
15'b0000101001011110011 : color = 12'he73;
15'b0000101001011110100 : color = 12'he73;
15'b0000101000100110011 : color = 12'he73;
15'b0000101000100110100 : color = 12'he73;
15'b0000101000100110101 : color = 12'he73;
15'b0000101000100110110 : color = 12'he73;
15'b0000101000100110111 : color = 12'he73;
15'b0000101000100111000 : color = 12'he73;
15'b0000101000100111001 : color = 12'he73;
15'b0000101000100111010 : color = 12'he73;
15'b0000101000100111011 : color = 12'he73;
15'b0000101000100111100 : color = 12'he73;
15'b0000101000100111101 : color = 12'he73;
15'b0000101000100111110 : color = 12'he73;
15'b0000101000100111111 : color = 12'he73;
15'b0000101000101000000 : color = 12'he61;
15'b0000101000101000001 : color = 12'hf00;
15'b0000101000101000010 : color = 12'hf01;
15'b0000101000101000011 : color = 12'hf73;
15'b0000101000101000100 : color = 12'he73;
15'b0000101000101000101 : color = 12'he73;
15'b0000101000101000110 : color = 12'he51;
15'b0000101000101000111 : color = 12'hf63;
15'b0000101000101001000 : color = 12'he73;
15'b0000101000101001001 : color = 12'he73;
15'b0000101000101001010 : color = 12'he73;
15'b0000101000101001011 : color = 12'he51;
15'b0000101000101001100 : color = 12'hf00;
15'b0000101000101001101 : color = 12'hf41;
15'b0000101000101001110 : color = 12'hf42;
15'b0000101000101001111 : color = 12'he73;
15'b0000101000101010000 : color = 12'he73;
15'b0000101000101010001 : color = 12'he73;
15'b0000101000101010010 : color = 12'he73;
15'b0000101000101010011 : color = 12'he73;
15'b0000101000101010100 : color = 12'he73;
15'b0000101000101010101 : color = 12'he73;
15'b0000101000101010110 : color = 12'he73;
15'b0000101000101010111 : color = 12'he73;
15'b0000101000101011000 : color = 12'he73;
15'b0000101000101011001 : color = 12'he73;
15'b0000101000101011010 : color = 12'he73;
15'b0000101000101011011 : color = 12'he73;
15'b0000101000101011100 : color = 12'he73;
15'b0000101000101011101 : color = 12'he73;
15'b0000101000101011110 : color = 12'he73;
15'b0000101000101011111 : color = 12'he73;
15'b0000101000101100000 : color = 12'he73;
15'b0000101000101100001 : color = 12'he73;
15'b0000101000101100010 : color = 12'he73;
15'b0000101000101100011 : color = 12'he73;
15'b0000101000101100100 : color = 12'he73;
15'b0000101000101100101 : color = 12'he73;
15'b0000101000101100110 : color = 12'he73;
15'b0000101000101100111 : color = 12'he73;
15'b0000101000101101000 : color = 12'he73;
15'b0000101000101101001 : color = 12'he73;
15'b0000101000101101010 : color = 12'he73;
15'b0000101000101101011 : color = 12'he51;
15'b0000101000101101100 : color = 12'hf00;
15'b0000101000101101101 : color = 12'hf63;
15'b0000101000101101110 : color = 12'he73;
15'b0000101000101101111 : color = 12'he73;
15'b0000101000101110000 : color = 12'he61;
15'b0000101000101110001 : color = 12'hf00;
15'b0000101000101110010 : color = 12'hf53;
15'b0000101000101110011 : color = 12'he73;
15'b0000101000101110100 : color = 12'he73;
15'b0000101000101110101 : color = 12'he73;
15'b0000101000101110110 : color = 12'he73;
15'b0000101000101110111 : color = 12'he72;
15'b0000101000101111000 : color = 12'hf10;
15'b0000101000101111001 : color = 12'hf32;
15'b0000101000101111010 : color = 12'he73;
15'b0000101000101111011 : color = 12'he73;
15'b0000101000101111100 : color = 12'he73;
15'b0000101000101111101 : color = 12'he72;
15'b0000101000101111110 : color = 12'hf10;
15'b0000101000101111111 : color = 12'hf32;
15'b0000101000110000000 : color = 12'he73;
15'b0000101000110000001 : color = 12'he73;
15'b0000101000110000010 : color = 12'he73;
15'b0000101000110000011 : color = 12'he73;
15'b0000101000110000100 : color = 12'he73;
15'b0000101000110000101 : color = 12'he73;
15'b0000101000110000110 : color = 12'he73;
15'b0000101000110000111 : color = 12'he73;
15'b0000101000110001000 : color = 12'he73;
15'b0000101000110001001 : color = 12'he73;
15'b0000101000110001010 : color = 12'he73;
15'b0000101000110001011 : color = 12'he73;
15'b0000101000110001100 : color = 12'he73;
15'b0000101000110001101 : color = 12'he73;
15'b0000101000110001110 : color = 12'he73;
15'b0000101000110001111 : color = 12'he73;
15'b0000101000110010000 : color = 12'he73;
15'b0000101000110010001 : color = 12'he73;
15'b0000101000110010010 : color = 12'he73;
15'b0000101000110010011 : color = 12'hf51;
15'b0000101000110010100 : color = 12'hf31;
15'b0000101000110010101 : color = 12'hf31;
15'b0000101000110010110 : color = 12'hf31;
15'b0000101000110010111 : color = 12'hf31;
15'b0000101000110011000 : color = 12'hf31;
15'b0000101000110011001 : color = 12'hf31;
15'b0000101000110011010 : color = 12'hf31;
15'b0000101000110011011 : color = 12'hf31;
15'b0000101000110011100 : color = 12'hf31;
15'b0000101000110011101 : color = 12'hf31;
15'b0000101000110011110 : color = 12'hf31;
15'b0000101000110011111 : color = 12'hf10;
15'b0000101000110100000 : color = 12'hf00;
15'b0000101000110100001 : color = 12'hf11;
15'b0000101000110100010 : color = 12'hf31;
15'b0000101000110100011 : color = 12'hf10;
15'b0000101000110100100 : color = 12'hf31;
15'b0000101000110100101 : color = 12'hf31;
15'b0000101000110100110 : color = 12'hf31;
15'b0000101000110100111 : color = 12'hf31;
15'b0000101000110101000 : color = 12'hf31;
15'b0000101000110101001 : color = 12'hf30;
15'b0000101000110101010 : color = 12'hf00;
15'b0000101000110101011 : color = 12'hf00;
15'b0000101000110101100 : color = 12'hf00;
15'b0000101000110101101 : color = 12'hf63;
15'b0000101000110101110 : color = 12'he73;
15'b0000101000110101111 : color = 12'he73;
15'b0000101000110110000 : color = 12'he73;
15'b0000101000110110001 : color = 12'he73;
15'b0000101000110110010 : color = 12'he73;
15'b0000101000110110011 : color = 12'he73;
15'b0000101000110110100 : color = 12'he73;
15'b0000101000110110101 : color = 12'he73;
15'b0000101000110110110 : color = 12'he73;
15'b0000101000110110111 : color = 12'he73;
15'b0000101000110111000 : color = 12'he73;
15'b0000101000110111001 : color = 12'he73;
15'b0000101000110111010 : color = 12'he73;
15'b0000101000110111011 : color = 12'he73;
15'b0000101000110111100 : color = 12'he73;
15'b0000101000110111101 : color = 12'he73;
15'b0000101000110111110 : color = 12'he73;
15'b0000101000110111111 : color = 12'he73;
15'b0000101000111000000 : color = 12'he73;
15'b0000101000111000001 : color = 12'he73;
15'b0000101000111000010 : color = 12'he73;
15'b0000101000111000011 : color = 12'he73;
15'b0000101000111000100 : color = 12'he73;
15'b0000101000111000101 : color = 12'he73;
15'b0000101000111000110 : color = 12'he72;
15'b0000101000111000111 : color = 12'hf00;
15'b0000101000111001000 : color = 12'hf42;
15'b0000101000111001001 : color = 12'he73;
15'b0000101000111001010 : color = 12'he73;
15'b0000101000111001011 : color = 12'he73;
15'b0000101000111001100 : color = 12'he73;
15'b0000101000111001101 : color = 12'he73;
15'b0000101000111001110 : color = 12'he73;
15'b0000101000111001111 : color = 12'he73;
15'b0000101000111010000 : color = 12'he72;
15'b0000101000111010001 : color = 12'hf10;
15'b0000101000111010010 : color = 12'hf32;
15'b0000101000111010011 : color = 12'he73;
15'b0000101000111010100 : color = 12'he73;
15'b0000101000111010101 : color = 12'he73;
15'b0000101000111010110 : color = 12'hf40;
15'b0000101000111010111 : color = 12'hf01;
15'b0000101000111011000 : color = 12'hf73;
15'b0000101000111011001 : color = 12'he73;
15'b0000101000111011010 : color = 12'he73;
15'b0000101000111011011 : color = 12'he73;
15'b0000101000111011100 : color = 12'he73;
15'b0000101000111011101 : color = 12'he73;
15'b0000101000111011110 : color = 12'he73;
15'b0000101000111011111 : color = 12'he73;
15'b0000101000111100000 : color = 12'he73;
15'b0000101000111100001 : color = 12'he73;
15'b0000101000111100010 : color = 12'he73;
15'b0000101000111100011 : color = 12'he73;
15'b0000101000111100100 : color = 12'he73;
15'b0000101000111100101 : color = 12'he73;
15'b0000101000111100110 : color = 12'he73;
15'b0000101000111100111 : color = 12'he73;
15'b0000101000111101000 : color = 12'he73;
15'b0000101000111101001 : color = 12'he73;
15'b0000101000111101010 : color = 12'he73;
15'b0000101000111101011 : color = 12'he73;
15'b0000101000111101100 : color = 12'he73;
15'b0000101000111101101 : color = 12'hf40;
15'b0000101000111101110 : color = 12'hf31;
15'b0000101000111101111 : color = 12'hf63;
15'b0000101000111110000 : color = 12'he73;
15'b0000101000111110001 : color = 12'he73;
15'b0000101000111110010 : color = 12'he73;
15'b0000101000111110011 : color = 12'he72;
15'b0000101000111110100 : color = 12'hf32;
15'b0000101000111110101 : color = 12'he73;
15'b0000101000111110110 : color = 12'he73;
15'b0000101000111110111 : color = 12'he73;
15'b0000101000111111000 : color = 12'he73;
15'b0000101000111111001 : color = 12'he73;
15'b0000101000111111010 : color = 12'he73;
15'b0000101000111111011 : color = 12'hf30;
15'b0000101000111111100 : color = 12'hf00;
15'b0000101000111111101 : color = 12'hf53;
15'b0000101000111111110 : color = 12'he73;
15'b0000101000111111111 : color = 12'he73;
15'b0000101001000000000 : color = 12'he73;
15'b0000101001000000001 : color = 12'he51;
15'b0000101001000000010 : color = 12'hf32;
15'b0000101001000000011 : color = 12'he73;
15'b0000101001000000100 : color = 12'he73;
15'b0000101001000000101 : color = 12'he73;
15'b0000101001000000110 : color = 12'he73;
15'b0000101001000000111 : color = 12'he73;
15'b0000101001000001000 : color = 12'he73;
15'b0000101001000001001 : color = 12'he73;
15'b0000101001000001010 : color = 12'he73;
15'b0000101001000001011 : color = 12'he73;
15'b0000101001000001100 : color = 12'he73;
15'b0000101001000001101 : color = 12'he73;
15'b0000101001000001110 : color = 12'he73;
15'b0000101001000001111 : color = 12'he73;
15'b0000101001000010000 : color = 12'he73;
15'b0000101001000010001 : color = 12'he73;
15'b0000101001000010010 : color = 12'he73;
15'b0000101001000010011 : color = 12'he73;
15'b0000101001000010100 : color = 12'he73;
15'b0000101001000010101 : color = 12'he73;
15'b0000101001000010110 : color = 12'he73;
15'b0000101001000010111 : color = 12'he73;
15'b0000101001000011000 : color = 12'he73;
15'b0000101001000011001 : color = 12'he73;
15'b0000101001000011010 : color = 12'he73;
15'b0000101001000011011 : color = 12'he51;
15'b0000101001000011100 : color = 12'hf00;
15'b0000101001000011101 : color = 12'hf63;
15'b0000101001000011110 : color = 12'he73;
15'b0000101001000011111 : color = 12'he73;
15'b0000101001000100000 : color = 12'hf40;
15'b0000101001000100001 : color = 12'hf11;
15'b0000101001000100010 : color = 12'hf73;
15'b0000101001000100011 : color = 12'he73;
15'b0000101001000100100 : color = 12'he73;
15'b0000101001000100101 : color = 12'he73;
15'b0000101001000100110 : color = 12'he61;
15'b0000101001000100111 : color = 12'hf00;
15'b0000101001000101000 : color = 12'hf53;
15'b0000101001000101001 : color = 12'he73;
15'b0000101001000101010 : color = 12'he73;
15'b0000101001000101011 : color = 12'he73;
15'b0000101001000101100 : color = 12'he73;
15'b0000101001000101101 : color = 12'he51;
15'b0000101001000101110 : color = 12'hf00;
15'b0000101001000101111 : color = 12'hf63;
15'b0000101001000110000 : color = 12'he73;
15'b0000101001000110001 : color = 12'he73;
15'b0000101001000110010 : color = 12'he73;
15'b0000101001000110011 : color = 12'he73;
15'b0000101001000110100 : color = 12'he73;
15'b0000101001000110101 : color = 12'he73;
15'b0000101001000110110 : color = 12'he73;
15'b0000101001000110111 : color = 12'he73;
15'b0000101001000111000 : color = 12'he73;
15'b0000101001000111001 : color = 12'he73;
15'b0000101001000111010 : color = 12'he73;
15'b0000101001000111011 : color = 12'he73;
15'b0000101001000111100 : color = 12'he73;
15'b0000101001000111101 : color = 12'he73;
15'b0000101001000111110 : color = 12'he73;
15'b0000101001000111111 : color = 12'he73;
15'b0000101001001000000 : color = 12'he73;
15'b0000101001001000001 : color = 12'he73;
15'b0000101001001000010 : color = 12'he73;
15'b0000101001001000011 : color = 12'he62;
15'b0000101001001000100 : color = 12'hf62;
15'b0000101001001000101 : color = 12'he73;
15'b0000101001001000110 : color = 12'he73;
15'b0000101001001000111 : color = 12'he73;
15'b0000101001001001000 : color = 12'hf40;
15'b0000101001001001001 : color = 12'hf01;
15'b0000101001001001010 : color = 12'hf73;
15'b0000101001001001011 : color = 12'he73;
15'b0000101001001001100 : color = 12'he73;
15'b0000101001001001101 : color = 12'he73;
15'b0000101001001001110 : color = 12'he73;
15'b0000101001001001111 : color = 12'he73;
15'b0000101001001010000 : color = 12'he73;
15'b0000101001001010001 : color = 12'he73;
15'b0000101001001010010 : color = 12'he73;
15'b0000101001001010011 : color = 12'he73;
15'b0000101001001010100 : color = 12'he51;
15'b0000101001001010101 : color = 12'hf00;
15'b0000101001001010110 : color = 12'hf53;
15'b0000101001001010111 : color = 12'he73;
15'b0000101001001011000 : color = 12'he73;
15'b0000101001001011001 : color = 12'he73;
15'b0000101001001011010 : color = 12'he73;
15'b0000101001001011011 : color = 12'he73;
15'b0000101001001011100 : color = 12'he73;
15'b0000101001001011101 : color = 12'he73;
15'b0000101001001011110 : color = 12'he73;
15'b0000101001001011111 : color = 12'he73;
15'b0000101001001100000 : color = 12'he73;
15'b0000101001001100001 : color = 12'he73;
15'b0000101001001100010 : color = 12'he73;
15'b0000101001001100011 : color = 12'he73;
15'b0000101001001100100 : color = 12'he73;
15'b0000101001001100101 : color = 12'he73;
15'b0000101001001100110 : color = 12'he73;
15'b0000101001001100111 : color = 12'he73;
15'b0000101001001101000 : color = 12'he73;
15'b0000101001001101001 : color = 12'he73;
15'b0000101001001101010 : color = 12'he73;
15'b0000101001001101011 : color = 12'he73;
15'b0000101001001101100 : color = 12'he73;
15'b0000101001001101101 : color = 12'he73;
15'b0000101001001101110 : color = 12'he73;
15'b0000101001001101111 : color = 12'he73;
15'b0000101001001110000 : color = 12'he73;
15'b0000101001001110001 : color = 12'he73;
15'b0000101001001110010 : color = 12'he73;
15'b0000101001001110011 : color = 12'he73;
15'b0000101001001110100 : color = 12'he73;
15'b0000101001001110101 : color = 12'hf30;
15'b0000101001001110110 : color = 12'hf11;
15'b0000101001001110111 : color = 12'hf73;
15'b0000101001001111000 : color = 12'he73;
15'b0000101001001111001 : color = 12'he73;
15'b0000101001001111010 : color = 12'he73;
15'b0000101001001111011 : color = 12'he73;
15'b0000101001001111100 : color = 12'he73;
15'b0000101001001111101 : color = 12'he73;
15'b0000101001001111110 : color = 12'he73;
15'b0000101001001111111 : color = 12'he73;
15'b0000101001010000000 : color = 12'he72;
15'b0000101001010000001 : color = 12'hf10;
15'b0000101001010000010 : color = 12'hf32;
15'b0000101001010000011 : color = 12'he73;
15'b0000101001010000100 : color = 12'he73;
15'b0000101001010000101 : color = 12'he73;
15'b0000101001010000110 : color = 12'he73;
15'b0000101001010000111 : color = 12'he73;
15'b0000101001010001000 : color = 12'he73;
15'b0000101001010001001 : color = 12'he73;
15'b0000101001010001010 : color = 12'he73;
15'b0000101001010001011 : color = 12'he73;
15'b0000101001010001100 : color = 12'he73;
15'b0000101001010001101 : color = 12'he73;
15'b0000101001010001110 : color = 12'he73;
15'b0000101001010001111 : color = 12'he73;
15'b0000101001010010000 : color = 12'he73;
15'b0000101001010010001 : color = 12'he73;
15'b0000101001010010010 : color = 12'he73;
15'b0000101001010010011 : color = 12'he73;
15'b0000101001010010100 : color = 12'he73;
15'b0000101001010010101 : color = 12'he73;
15'b0000101001010010110 : color = 12'he73;
15'b0000101001010010111 : color = 12'he73;
15'b0000101001010011000 : color = 12'he73;
15'b0000101001010011001 : color = 12'he73;
15'b0000101001010011010 : color = 12'he73;
15'b0000101001010011011 : color = 12'he73;
15'b0000101001010011100 : color = 12'he72;
15'b0000101001010011101 : color = 12'hf63;
15'b0000101001010011110 : color = 12'he73;
15'b0000101001010011111 : color = 12'he72;
15'b0000101001010100000 : color = 12'hf10;
15'b0000101001010100001 : color = 12'hf32;
15'b0000101001010100010 : color = 12'he73;
15'b0000101001010100011 : color = 12'he73;
15'b0000101001010100100 : color = 12'he73;
15'b0000101001010100101 : color = 12'he73;
15'b0000101001010100110 : color = 12'he51;
15'b0000101001010100111 : color = 12'hf00;
15'b0000101001010101000 : color = 12'hf31;
15'b0000101001010101001 : color = 12'hf31;
15'b0000101001010101010 : color = 12'hf31;
15'b0000101001010101011 : color = 12'hf31;
15'b0000101001010101100 : color = 12'hf10;
15'b0000101001010101101 : color = 12'hf10;
15'b0000101001010101110 : color = 12'hf31;
15'b0000101001010101111 : color = 12'hf31;
15'b0000101001010110000 : color = 12'hf31;
15'b0000101001010110001 : color = 12'hf30;
15'b0000101001010110010 : color = 12'hf00;
15'b0000101001010110011 : color = 12'hf63;
15'b0000101001010110100 : color = 12'he73;
15'b0000101001010110101 : color = 12'he73;
15'b0000101001010110110 : color = 12'he73;
15'b0000101001010110111 : color = 12'he73;
15'b0000101001010111000 : color = 12'he73;
15'b0000101001010111001 : color = 12'he73;
15'b0000101001010111010 : color = 12'he73;
15'b0000101001010111011 : color = 12'he73;
15'b0000101001010111100 : color = 12'he73;
15'b0000101001010111101 : color = 12'he73;
15'b0000101001010111110 : color = 12'he73;
15'b0000101001010111111 : color = 12'he73;
15'b0000101001011000000 : color = 12'he73;
15'b0000101001011000001 : color = 12'he73;
15'b0000101001011000010 : color = 12'he73;
15'b0000101001011000011 : color = 12'he73;
15'b0000101001011000100 : color = 12'he73;
15'b0000101001011000101 : color = 12'he73;
15'b0000101001011000110 : color = 12'he73;
15'b0000101001011000111 : color = 12'he73;
15'b0000101001011001000 : color = 12'he73;
15'b0000101001011001001 : color = 12'he73;
15'b0000101001011001010 : color = 12'he73;
15'b0000101001011001011 : color = 12'he73;
15'b0000101001011001100 : color = 12'he73;
15'b0000101001011001101 : color = 12'he73;
15'b0000101001011001110 : color = 12'he73;
15'b0000101001011001111 : color = 12'he62;
15'b0000101001011010000 : color = 12'hf10;
15'b0000101001011010001 : color = 12'hf11;
15'b0000101001011010010 : color = 12'hf52;
15'b0000101001011010011 : color = 12'he73;
15'b0000101001011010100 : color = 12'he73;
15'b0000101001011010101 : color = 12'he73;
15'b0000101001011010110 : color = 12'he73;
15'b0000101001011010111 : color = 12'he73;
15'b0000101001011011000 : color = 12'he73;
15'b0000101001011011001 : color = 12'he73;
15'b0000101001011011010 : color = 12'he61;
15'b0000101001011011011 : color = 12'hf00;
15'b0000101001011011100 : color = 12'hf00;
15'b0000101001011011101 : color = 12'hf52;
15'b0000101001011011110 : color = 12'he73;
15'b0000101001011011111 : color = 12'he73;
15'b0000101001011100000 : color = 12'he73;
15'b0000101001011100001 : color = 12'he73;
15'b0000101001011100010 : color = 12'he73;
15'b0000101001011100011 : color = 12'he73;
15'b0000101001011100100 : color = 12'he73;
15'b0000101001011100101 : color = 12'he73;
15'b0000101001011100110 : color = 12'he73;
15'b0000101001011100111 : color = 12'he73;
15'b0000101001011101000 : color = 12'he73;
15'b0000101001011101001 : color = 12'he73;
15'b0000101001011101010 : color = 12'he73;
15'b0000101001011101011 : color = 12'he73;
15'b0000101001011101100 : color = 12'he73;
15'b0000101001011101101 : color = 12'he73;
15'b0000101001011101110 : color = 12'he73;
15'b0000101001011101111 : color = 12'he73;
15'b0000101001011110000 : color = 12'he73;
15'b0000101001011110001 : color = 12'he73;
15'b0000101001011110010 : color = 12'he73;
15'b0000101001011110011 : color = 12'he73;
15'b0000101001011110100 : color = 12'he73;
15'b0000101001011110101 : color = 12'he73;
15'b0000101001011110110 : color = 12'he72;
15'b0000101001011110111 : color = 12'hf10;
15'b0000101001011111000 : color = 12'hf42;
15'b0000101001011111001 : color = 12'he73;
15'b0000101001011111010 : color = 12'he73;
15'b0000101001011111011 : color = 12'he73;
15'b0000101001011111100 : color = 12'he73;
15'b0000101001011111101 : color = 12'he73;
15'b0000101001011111110 : color = 12'he61;
15'b0000101001011111111 : color = 12'hf10;
15'b0000101001100000000 : color = 12'hf52;
15'b0000101001100000001 : color = 12'hf73;
15'b0000101001100000010 : color = 12'he62;
15'b0000101001100000011 : color = 12'hf63;
15'b0000101001100000100 : color = 12'he73;
15'b0000101001100000101 : color = 12'he73;
15'b0000101001100000110 : color = 12'hf30;
15'b0000101001100000111 : color = 12'hf11;
15'b0000101001100001000 : color = 12'hf73;
15'b0000101001100001001 : color = 12'he73;
15'b0000101001100001010 : color = 12'he72;
15'b0000101001100001011 : color = 12'hf11;
15'b0000101001100001100 : color = 12'hf73;
15'b0000101001100001101 : color = 12'he73;
15'b0000101001100001110 : color = 12'he73;
15'b0000101001100001111 : color = 12'he73;
15'b0000101001100010000 : color = 12'he73;
15'b0000101001100010001 : color = 12'he73;
15'b0000101001100010010 : color = 12'he73;
15'b0000101001100010011 : color = 12'he73;
15'b0000101001100010100 : color = 12'he73;
15'b0000101001100010101 : color = 12'he73;
15'b0000101001100010110 : color = 12'he73;
15'b0000101001100010111 : color = 12'he73;
15'b0000101001100011000 : color = 12'he73;
15'b0000101001100011001 : color = 12'he73;
15'b0000101001100011010 : color = 12'he73;
15'b0000101001100011011 : color = 12'he73;
15'b0000101001100011100 : color = 12'he73;
15'b0000101001100011101 : color = 12'he73;
15'b0000101000101011100 : color = 12'he73;
15'b0000101000101011101 : color = 12'he73;
15'b0000101000101011110 : color = 12'he73;
15'b0000101000101011111 : color = 12'he73;
15'b0000101000101100000 : color = 12'he73;
15'b0000101000101100001 : color = 12'he73;
15'b0000101000101100010 : color = 12'he73;
15'b0000101000101100011 : color = 12'he73;
15'b0000101000101100100 : color = 12'he73;
15'b0000101000101100101 : color = 12'he73;
15'b0000101000101100110 : color = 12'he73;
15'b0000101000101100111 : color = 12'he73;
15'b0000101000101101000 : color = 12'he73;
15'b0000101000101101001 : color = 12'he72;
15'b0000101000101101010 : color = 12'hf00;
15'b0000101000101101011 : color = 12'hf00;
15'b0000101000101101100 : color = 12'hf53;
15'b0000101000101101101 : color = 12'he73;
15'b0000101000101101110 : color = 12'he73;
15'b0000101000101101111 : color = 12'he73;
15'b0000101000101110000 : color = 12'he73;
15'b0000101000101110001 : color = 12'he73;
15'b0000101000101110010 : color = 12'he73;
15'b0000101000101110011 : color = 12'he73;
15'b0000101000101110100 : color = 12'hf40;
15'b0000101000101110101 : color = 12'hf01;
15'b0000101000101110110 : color = 12'hf61;
15'b0000101000101110111 : color = 12'hf32;
15'b0000101000101111000 : color = 12'he73;
15'b0000101000101111001 : color = 12'he73;
15'b0000101000101111010 : color = 12'he73;
15'b0000101000101111011 : color = 12'he73;
15'b0000101000101111100 : color = 12'he73;
15'b0000101000101111101 : color = 12'he73;
15'b0000101000101111110 : color = 12'he73;
15'b0000101000101111111 : color = 12'he73;
15'b0000101000110000000 : color = 12'he73;
15'b0000101000110000001 : color = 12'he73;
15'b0000101000110000010 : color = 12'he73;
15'b0000101000110000011 : color = 12'he73;
15'b0000101000110000100 : color = 12'he73;
15'b0000101000110000101 : color = 12'he73;
15'b0000101000110000110 : color = 12'he73;
15'b0000101000110000111 : color = 12'he73;
15'b0000101000110001000 : color = 12'he73;
15'b0000101000110001001 : color = 12'he73;
15'b0000101000110001010 : color = 12'he73;
15'b0000101000110001011 : color = 12'he73;
15'b0000101000110001100 : color = 12'he73;
15'b0000101000110001101 : color = 12'he73;
15'b0000101000110001110 : color = 12'he73;
15'b0000101000110001111 : color = 12'he73;
15'b0000101000110010000 : color = 12'he73;
15'b0000101000110010001 : color = 12'he73;
15'b0000101000110010010 : color = 12'he73;
15'b0000101000110010011 : color = 12'he73;
15'b0000101000110010100 : color = 12'he51;
15'b0000101000110010101 : color = 12'hf00;
15'b0000101000110010110 : color = 12'hf63;
15'b0000101000110010111 : color = 12'he73;
15'b0000101000110011000 : color = 12'he73;
15'b0000101000110011001 : color = 12'he61;
15'b0000101000110011010 : color = 12'hf00;
15'b0000101000110011011 : color = 12'hf53;
15'b0000101000110011100 : color = 12'he73;
15'b0000101000110011101 : color = 12'he73;
15'b0000101000110011110 : color = 12'he73;
15'b0000101000110011111 : color = 12'hf52;
15'b0000101000110100000 : color = 12'hf62;
15'b0000101000110100001 : color = 12'hf10;
15'b0000101000110100010 : color = 12'hf32;
15'b0000101000110100011 : color = 12'he73;
15'b0000101000110100100 : color = 12'he73;
15'b0000101000110100101 : color = 12'he73;
15'b0000101000110100110 : color = 12'he72;
15'b0000101000110100111 : color = 12'hf10;
15'b0000101000110101000 : color = 12'hf32;
15'b0000101000110101001 : color = 12'he73;
15'b0000101000110101010 : color = 12'he73;
15'b0000101000110101011 : color = 12'he73;
15'b0000101000110101100 : color = 12'he73;
15'b0000101000110101101 : color = 12'he73;
15'b0000101000110101110 : color = 12'he73;
15'b0000101000110101111 : color = 12'he73;
15'b0000101000110110000 : color = 12'he73;
15'b0000101000110110001 : color = 12'he73;
15'b0000101000110110010 : color = 12'he73;
15'b0000101000110110011 : color = 12'he73;
15'b0000101000110110100 : color = 12'he73;
15'b0000101000110110101 : color = 12'he73;
15'b0000101000110110110 : color = 12'he73;
15'b0000101000110110111 : color = 12'he73;
15'b0000101000110111000 : color = 12'he73;
15'b0000101000110111001 : color = 12'he73;
15'b0000101000110111010 : color = 12'he73;
15'b0000101000110111011 : color = 12'he73;
15'b0000101000110111100 : color = 12'he73;
15'b0000101000110111101 : color = 12'hf62;
15'b0000101000110111110 : color = 12'hf73;
15'b0000101000110111111 : color = 12'he73;
15'b0000101000111000000 : color = 12'he73;
15'b0000101000111000001 : color = 12'he73;
15'b0000101000111000010 : color = 12'he73;
15'b0000101000111000011 : color = 12'he73;
15'b0000101000111000100 : color = 12'he73;
15'b0000101000111000101 : color = 12'he73;
15'b0000101000111000110 : color = 12'he72;
15'b0000101000111000111 : color = 12'hf00;
15'b0000101000111001000 : color = 12'hf00;
15'b0000101000111001001 : color = 12'hf00;
15'b0000101000111001010 : color = 12'hf52;
15'b0000101000111001011 : color = 12'hf32;
15'b0000101000111001100 : color = 12'he73;
15'b0000101000111001101 : color = 12'he73;
15'b0000101000111001110 : color = 12'he73;
15'b0000101000111001111 : color = 12'he73;
15'b0000101000111010000 : color = 12'he73;
15'b0000101000111010001 : color = 12'he73;
15'b0000101000111010010 : color = 12'he73;
15'b0000101000111010011 : color = 12'he73;
15'b0000101000111010100 : color = 12'he73;
15'b0000101000111010101 : color = 12'he73;
15'b0000101000111010110 : color = 12'he73;
15'b0000101000111010111 : color = 12'he73;
15'b0000101000111011000 : color = 12'he73;
15'b0000101000111011001 : color = 12'he73;
15'b0000101000111011010 : color = 12'he73;
15'b0000101000111011011 : color = 12'he73;
15'b0000101000111011100 : color = 12'he73;
15'b0000101000111011101 : color = 12'he73;
15'b0000101000111011110 : color = 12'he73;
15'b0000101000111011111 : color = 12'he73;
15'b0000101000111100000 : color = 12'he73;
15'b0000101000111100001 : color = 12'he73;
15'b0000101000111100010 : color = 12'he73;
15'b0000101000111100011 : color = 12'he73;
15'b0000101000111100100 : color = 12'he73;
15'b0000101000111100101 : color = 12'he73;
15'b0000101000111100110 : color = 12'he73;
15'b0000101000111100111 : color = 12'he73;
15'b0000101000111101000 : color = 12'he73;
15'b0000101000111101001 : color = 12'he73;
15'b0000101000111101010 : color = 12'he73;
15'b0000101000111101011 : color = 12'he73;
15'b0000101000111101100 : color = 12'he73;
15'b0000101000111101101 : color = 12'he73;
15'b0000101000111101110 : color = 12'he73;
15'b0000101000111101111 : color = 12'he72;
15'b0000101000111110000 : color = 12'hf00;
15'b0000101000111110001 : color = 12'hf42;
15'b0000101000111110010 : color = 12'he73;
15'b0000101000111110011 : color = 12'he73;
15'b0000101000111110100 : color = 12'he73;
15'b0000101000111110101 : color = 12'he73;
15'b0000101000111110110 : color = 12'he73;
15'b0000101000111110111 : color = 12'he73;
15'b0000101000111111000 : color = 12'he73;
15'b0000101000111111001 : color = 12'he72;
15'b0000101000111111010 : color = 12'hf10;
15'b0000101000111111011 : color = 12'hf32;
15'b0000101000111111100 : color = 12'he73;
15'b0000101000111111101 : color = 12'he73;
15'b0000101000111111110 : color = 12'he73;
15'b0000101000111111111 : color = 12'hf40;
15'b0000101001000000000 : color = 12'hf01;
15'b0000101001000000001 : color = 12'hf73;
15'b0000101001000000010 : color = 12'he73;
15'b0000101001000000011 : color = 12'he73;
15'b0000101001000000100 : color = 12'he73;
15'b0000101001000000101 : color = 12'he73;
15'b0000101001000000110 : color = 12'he73;
15'b0000101001000000111 : color = 12'he73;
15'b0000101001000001000 : color = 12'he73;
15'b0000101001000001001 : color = 12'he73;
15'b0000101001000001010 : color = 12'he73;
15'b0000101001000001011 : color = 12'he73;
15'b0000101001000001100 : color = 12'he73;
15'b0000101001000001101 : color = 12'he73;
15'b0000101001000001110 : color = 12'he73;
15'b0000101001000001111 : color = 12'he73;
15'b0000101001000010000 : color = 12'he73;
15'b0000101001000010001 : color = 12'he73;
15'b0000101001000010010 : color = 12'he73;
15'b0000101001000010011 : color = 12'he73;
15'b0000101001000010100 : color = 12'he72;
15'b0000101001000010101 : color = 12'hf41;
15'b0000101001000010110 : color = 12'hf63;
15'b0000101001000010111 : color = 12'he73;
15'b0000101001000011000 : color = 12'he73;
15'b0000101001000011001 : color = 12'he73;
15'b0000101001000011010 : color = 12'he73;
15'b0000101001000011011 : color = 12'he73;
15'b0000101001000011100 : color = 12'he73;
15'b0000101001000011101 : color = 12'hf30;
15'b0000101001000011110 : color = 12'hf63;
15'b0000101001000011111 : color = 12'he73;
15'b0000101001000100000 : color = 12'he73;
15'b0000101001000100001 : color = 12'he73;
15'b0000101001000100010 : color = 12'he73;
15'b0000101001000100011 : color = 12'he61;
15'b0000101001000100100 : color = 12'hf00;
15'b0000101001000100101 : color = 12'hf11;
15'b0000101001000100110 : color = 12'hf73;
15'b0000101001000100111 : color = 12'he73;
15'b0000101001000101000 : color = 12'he73;
15'b0000101001000101001 : color = 12'he73;
15'b0000101001000101010 : color = 12'he73;
15'b0000101001000101011 : color = 12'he73;
15'b0000101001000101100 : color = 12'he73;
15'b0000101001000101101 : color = 12'he73;
15'b0000101001000101110 : color = 12'he73;
15'b0000101001000101111 : color = 12'he73;
15'b0000101001000110000 : color = 12'he73;
15'b0000101001000110001 : color = 12'he73;
15'b0000101001000110010 : color = 12'he73;
15'b0000101001000110011 : color = 12'he73;
15'b0000101001000110100 : color = 12'he73;
15'b0000101001000110101 : color = 12'he73;
15'b0000101001000110110 : color = 12'he73;
15'b0000101001000110111 : color = 12'he73;
15'b0000101001000111000 : color = 12'he73;
15'b0000101001000111001 : color = 12'he73;
15'b0000101001000111010 : color = 12'he73;
15'b0000101001000111011 : color = 12'he73;
15'b0000101001000111100 : color = 12'he73;
15'b0000101001000111101 : color = 12'he73;
15'b0000101001000111110 : color = 12'he73;
15'b0000101001000111111 : color = 12'he73;
15'b0000101001001000000 : color = 12'he73;
15'b0000101001001000001 : color = 12'he73;
15'b0000101001001000010 : color = 12'he73;
15'b0000101001001000011 : color = 12'he73;
15'b0000101001001000100 : color = 12'he51;
15'b0000101001001000101 : color = 12'hf00;
15'b0000101001001000110 : color = 12'hf63;
15'b0000101001001000111 : color = 12'he73;
15'b0000101001001001000 : color = 12'he73;
15'b0000101001001001001 : color = 12'hf40;
15'b0000101001001001010 : color = 12'hf11;
15'b0000101001001001011 : color = 12'hf73;
15'b0000101001001001100 : color = 12'he73;
15'b0000101001001001101 : color = 12'he73;
15'b0000101001001001110 : color = 12'he73;
15'b0000101001001001111 : color = 12'he61;
15'b0000101001001010000 : color = 12'hf00;
15'b0000101001001010001 : color = 12'hf53;
15'b0000101001001010010 : color = 12'he73;
15'b0000101001001010011 : color = 12'he73;
15'b0000101001001010100 : color = 12'he73;
15'b0000101001001010101 : color = 12'he73;
15'b0000101001001010110 : color = 12'he51;
15'b0000101001001010111 : color = 12'hf00;
15'b0000101001001011000 : color = 12'hf63;
15'b0000101001001011001 : color = 12'he73;
15'b0000101001001011010 : color = 12'he73;
15'b0000101001001011011 : color = 12'he73;
15'b0000101001001011100 : color = 12'he73;
15'b0000101001001011101 : color = 12'he73;
15'b0000101001001011110 : color = 12'he73;
15'b0000101001001011111 : color = 12'he73;
15'b0000101001001100000 : color = 12'he73;
15'b0000101001001100001 : color = 12'he73;
15'b0000101001001100010 : color = 12'he73;
15'b0000101001001100011 : color = 12'he73;
15'b0000101001001100100 : color = 12'he73;
15'b0000101001001100101 : color = 12'he73;
15'b0000101001001100110 : color = 12'he73;
15'b0000101001001100111 : color = 12'he73;
15'b0000101001001101000 : color = 12'he73;
15'b0000101001001101001 : color = 12'he73;
15'b0000101001001101010 : color = 12'he73;
15'b0000101001001101011 : color = 12'he73;
15'b0000101001001101100 : color = 12'he73;
15'b0000101001001101101 : color = 12'he73;
15'b0000101001001101110 : color = 12'he73;
15'b0000101001001101111 : color = 12'he73;
15'b0000101001001110000 : color = 12'he73;
15'b0000101001001110001 : color = 12'hf40;
15'b0000101001001110010 : color = 12'hf11;
15'b0000101001001110011 : color = 12'hf73;
15'b0000101001001110100 : color = 12'he73;
15'b0000101001001110101 : color = 12'he73;
15'b0000101001001110110 : color = 12'he73;
15'b0000101001001110111 : color = 12'he73;
15'b0000101001001111000 : color = 12'he73;
15'b0000101001001111001 : color = 12'he73;
15'b0000101001001111010 : color = 12'he73;
15'b0000101001001111011 : color = 12'he73;
15'b0000101001001111100 : color = 12'he73;
15'b0000101001001111101 : color = 12'he51;
15'b0000101001001111110 : color = 12'hf00;
15'b0000101001001111111 : color = 12'hf53;
15'b0000101001010000000 : color = 12'he73;
15'b0000101001010000001 : color = 12'he73;
15'b0000101001010000010 : color = 12'he73;
15'b0000101001010000011 : color = 12'he73;
15'b0000101001010000100 : color = 12'he73;
15'b0000101001010000101 : color = 12'he73;
15'b0000101001010000110 : color = 12'he73;
15'b0000101001010000111 : color = 12'he73;
15'b0000101001010001000 : color = 12'he73;
15'b0000101001010001001 : color = 12'he73;
15'b0000101001010001010 : color = 12'he73;
15'b0000101001010001011 : color = 12'he73;
15'b0000101001010001100 : color = 12'he73;
15'b0000101001010001101 : color = 12'he73;
15'b0000101001010001110 : color = 12'he73;
15'b0000101001010001111 : color = 12'he73;
15'b0000101001010010000 : color = 12'he73;
15'b0000101001010010001 : color = 12'he73;
15'b0000101001010010010 : color = 12'he73;
15'b0000101001010010011 : color = 12'he73;
15'b0000101001010010100 : color = 12'he73;
15'b0000101001010010101 : color = 12'he73;
15'b0000101001010010110 : color = 12'he73;
15'b0000101001010010111 : color = 12'he73;
15'b0000101001010011000 : color = 12'he73;
15'b0000101001010011001 : color = 12'he73;
15'b0000101001010011010 : color = 12'he73;
15'b0000101001010011011 : color = 12'he73;
15'b0000101001010011100 : color = 12'he73;
15'b0000101001010011101 : color = 12'he73;
15'b0000101001010011110 : color = 12'hf30;
15'b0000101001010011111 : color = 12'hf11;
15'b0000101001010100000 : color = 12'hf73;
15'b0000101001010100001 : color = 12'he73;
15'b0000101001010100010 : color = 12'he73;
15'b0000101001010100011 : color = 12'he73;
15'b0000101001010100100 : color = 12'he73;
15'b0000101001010100101 : color = 12'he73;
15'b0000101001010100110 : color = 12'he73;
15'b0000101001010100111 : color = 12'he73;
15'b0000101001010101000 : color = 12'he73;
15'b0000101001010101001 : color = 12'he72;
15'b0000101001010101010 : color = 12'hf10;
15'b0000101001010101011 : color = 12'hf32;
15'b0000101001010101100 : color = 12'he73;
15'b0000101001010101101 : color = 12'he73;
15'b0000101001010101110 : color = 12'he73;
15'b0000101001010101111 : color = 12'he73;
15'b0000101001010110000 : color = 12'he73;
15'b0000101001010110001 : color = 12'he73;
15'b0000101001010110010 : color = 12'he73;
15'b0000101001010110011 : color = 12'he73;
15'b0000101001010110100 : color = 12'he73;
15'b0000101001010110101 : color = 12'he73;
15'b0000101001010110110 : color = 12'he73;
15'b0000101001010110111 : color = 12'he73;
15'b0000101001010111000 : color = 12'he73;
15'b0000101001010111001 : color = 12'he73;
15'b0000101001010111010 : color = 12'he73;
15'b0000101001010111011 : color = 12'he73;
15'b0000101001010111100 : color = 12'he73;
15'b0000101001010111101 : color = 12'he73;
15'b0000101001010111110 : color = 12'he73;
15'b0000101001010111111 : color = 12'he73;
15'b0000101001011000000 : color = 12'he73;
15'b0000101001011000001 : color = 12'he73;
15'b0000101001011000010 : color = 12'he73;
15'b0000101001011000011 : color = 12'he73;
15'b0000101001011000100 : color = 12'he73;
15'b0000101001011000101 : color = 12'he73;
15'b0000101001011000110 : color = 12'he73;
15'b0000101001011000111 : color = 12'he73;
15'b0000101001011001000 : color = 12'he72;
15'b0000101001011001001 : color = 12'hf10;
15'b0000101001011001010 : color = 12'hf32;
15'b0000101001011001011 : color = 12'he73;
15'b0000101001011001100 : color = 12'he73;
15'b0000101001011001101 : color = 12'he73;
15'b0000101001011001110 : color = 12'he73;
15'b0000101001011001111 : color = 12'he51;
15'b0000101001011010000 : color = 12'hf00;
15'b0000101001011010001 : color = 12'hf63;
15'b0000101001011010010 : color = 12'he73;
15'b0000101001011010011 : color = 12'he73;
15'b0000101001011010100 : color = 12'he73;
15'b0000101001011010101 : color = 12'hf30;
15'b0000101001011010110 : color = 12'hf32;
15'b0000101001011010111 : color = 12'he73;
15'b0000101001011011000 : color = 12'he73;
15'b0000101001011011001 : color = 12'he73;
15'b0000101001011011010 : color = 12'he61;
15'b0000101001011011011 : color = 12'hf00;
15'b0000101001011011100 : color = 12'hf63;
15'b0000101001011011101 : color = 12'he73;
15'b0000101001011011110 : color = 12'he73;
15'b0000101001011011111 : color = 12'he73;
15'b0000101001011100000 : color = 12'he73;
15'b0000101001011100001 : color = 12'he73;
15'b0000101001011100010 : color = 12'he73;
15'b0000101001011100011 : color = 12'he73;
15'b0000101001011100100 : color = 12'he73;
15'b0000101001011100101 : color = 12'he73;
15'b0000101001011100110 : color = 12'he73;
15'b0000101001011100111 : color = 12'he73;
15'b0000101001011101000 : color = 12'he73;
15'b0000101001011101001 : color = 12'he73;
15'b0000101001011101010 : color = 12'he73;
15'b0000101001011101011 : color = 12'he73;
15'b0000101001011101100 : color = 12'he73;
15'b0000101001011101101 : color = 12'he73;
15'b0000101001011101110 : color = 12'he73;
15'b0000101001011101111 : color = 12'he73;
15'b0000101001011110000 : color = 12'he73;
15'b0000101001011110001 : color = 12'he73;
15'b0000101001011110010 : color = 12'he73;
15'b0000101001011110011 : color = 12'he73;
15'b0000101001011110100 : color = 12'he73;
15'b0000101001011110101 : color = 12'he73;
15'b0000101001011110110 : color = 12'hf62;
15'b0000101001011110111 : color = 12'hf10;
15'b0000101001011111000 : color = 12'hf00;
15'b0000101001011111001 : color = 12'hf52;
15'b0000101001011111010 : color = 12'hf73;
15'b0000101001011111011 : color = 12'he73;
15'b0000101001011111100 : color = 12'he73;
15'b0000101001011111101 : color = 12'he73;
15'b0000101001011111110 : color = 12'he73;
15'b0000101001011111111 : color = 12'he73;
15'b0000101001100000000 : color = 12'he73;
15'b0000101001100000001 : color = 12'he72;
15'b0000101001100000010 : color = 12'hf62;
15'b0000101001100000011 : color = 12'hf62;
15'b0000101001100000100 : color = 12'hf51;
15'b0000101001100000101 : color = 12'hf00;
15'b0000101001100000110 : color = 12'hf00;
15'b0000101001100000111 : color = 12'hf11;
15'b0000101001100001000 : color = 12'hf73;
15'b0000101001100001001 : color = 12'he73;
15'b0000101001100001010 : color = 12'he73;
15'b0000101001100001011 : color = 12'he73;
15'b0000101001100001100 : color = 12'he73;
15'b0000101001100001101 : color = 12'he73;
15'b0000101001100001110 : color = 12'he73;
15'b0000101001100001111 : color = 12'he73;
15'b0000101001100010000 : color = 12'he73;
15'b0000101001100010001 : color = 12'he73;
15'b0000101001100010010 : color = 12'he73;
15'b0000101001100010011 : color = 12'he73;
15'b0000101001100010100 : color = 12'he73;
15'b0000101001100010101 : color = 12'he73;
15'b0000101001100010110 : color = 12'he73;
15'b0000101001100010111 : color = 12'he73;
15'b0000101001100011000 : color = 12'he73;
15'b0000101001100011001 : color = 12'he73;
15'b0000101001100011010 : color = 12'he73;
15'b0000101001100011011 : color = 12'he73;
15'b0000101001100011100 : color = 12'he73;
15'b0000101001100011101 : color = 12'he73;
15'b0000101001100011110 : color = 12'he72;
15'b0000101001100011111 : color = 12'hf10;
15'b0000101001100100000 : color = 12'hf32;
15'b0000101001100100001 : color = 12'he73;
15'b0000101001100100010 : color = 12'he73;
15'b0000101001100100011 : color = 12'he73;
15'b0000101001100100100 : color = 12'he73;
15'b0000101001100100101 : color = 12'he73;
15'b0000101001100100110 : color = 12'he73;
15'b0000101001100100111 : color = 12'he73;
15'b0000101001100101000 : color = 12'he73;
15'b0000101001100101001 : color = 12'he73;
15'b0000101001100101010 : color = 12'he61;
15'b0000101001100101011 : color = 12'hf00;
15'b0000101001100101100 : color = 12'hf42;
15'b0000101001100101101 : color = 12'he73;
15'b0000101001100101110 : color = 12'he73;
15'b0000101001100101111 : color = 12'hf30;
15'b0000101001100110000 : color = 12'hf11;
15'b0000101001100110001 : color = 12'hf73;
15'b0000101001100110010 : color = 12'he73;
15'b0000101001100110011 : color = 12'he73;
15'b0000101001100110100 : color = 12'he73;
15'b0000101001100110101 : color = 12'he73;
15'b0000101001100110110 : color = 12'he73;
15'b0000101001100110111 : color = 12'he73;
15'b0000101001100111000 : color = 12'he73;
15'b0000101001100111001 : color = 12'he73;
15'b0000101001100111010 : color = 12'he73;
15'b0000101001100111011 : color = 12'he73;
15'b0000101001100111100 : color = 12'he73;
15'b0000101001100111101 : color = 12'he73;
15'b0000101001100111110 : color = 12'he73;
15'b0000101001100111111 : color = 12'he73;
15'b0000101001101000000 : color = 12'he73;
15'b0000101001101000001 : color = 12'he73;
15'b0000101001101000010 : color = 12'he73;
15'b0000101001101000011 : color = 12'he73;
15'b0000101001101000100 : color = 12'he73;
15'b0000101001101000101 : color = 12'he73;
15'b0000101001101000110 : color = 12'he73;
15'b0000101000110000101 : color = 12'he73;
15'b0000101000110000110 : color = 12'he73;
15'b0000101000110000111 : color = 12'he73;
15'b0000101000110001000 : color = 12'he73;
15'b0000101000110001001 : color = 12'he73;
15'b0000101000110001010 : color = 12'he73;
15'b0000101000110001011 : color = 12'he73;
15'b0000101000110001100 : color = 12'he73;
15'b0000101000110001101 : color = 12'he73;
15'b0000101000110001110 : color = 12'he73;
15'b0000101000110001111 : color = 12'he73;
15'b0000101000110010000 : color = 12'he73;
15'b0000101000110010001 : color = 12'he73;
15'b0000101000110010010 : color = 12'hf40;
15'b0000101000110010011 : color = 12'hf00;
15'b0000101000110010100 : color = 12'hf10;
15'b0000101000110010101 : color = 12'hf00;
15'b0000101000110010110 : color = 12'hf63;
15'b0000101000110010111 : color = 12'he73;
15'b0000101000110011000 : color = 12'he73;
15'b0000101000110011001 : color = 12'he73;
15'b0000101000110011010 : color = 12'he73;
15'b0000101000110011011 : color = 12'he73;
15'b0000101000110011100 : color = 12'he72;
15'b0000101000110011101 : color = 12'hf10;
15'b0000101000110011110 : color = 12'hf32;
15'b0000101000110011111 : color = 12'he72;
15'b0000101000110100000 : color = 12'hf01;
15'b0000101000110100001 : color = 12'hf73;
15'b0000101000110100010 : color = 12'he73;
15'b0000101000110100011 : color = 12'he73;
15'b0000101000110100100 : color = 12'he73;
15'b0000101000110100101 : color = 12'he73;
15'b0000101000110100110 : color = 12'he73;
15'b0000101000110100111 : color = 12'he73;
15'b0000101000110101000 : color = 12'he73;
15'b0000101000110101001 : color = 12'he73;
15'b0000101000110101010 : color = 12'he73;
15'b0000101000110101011 : color = 12'he73;
15'b0000101000110101100 : color = 12'he73;
15'b0000101000110101101 : color = 12'he73;
15'b0000101000110101110 : color = 12'he73;
15'b0000101000110101111 : color = 12'he73;
15'b0000101000110110000 : color = 12'he73;
15'b0000101000110110001 : color = 12'he73;
15'b0000101000110110010 : color = 12'he73;
15'b0000101000110110011 : color = 12'he73;
15'b0000101000110110100 : color = 12'he73;
15'b0000101000110110101 : color = 12'he73;
15'b0000101000110110110 : color = 12'he73;
15'b0000101000110110111 : color = 12'he73;
15'b0000101000110111000 : color = 12'he73;
15'b0000101000110111001 : color = 12'he73;
15'b0000101000110111010 : color = 12'he73;
15'b0000101000110111011 : color = 12'he73;
15'b0000101000110111100 : color = 12'he73;
15'b0000101000110111101 : color = 12'he51;
15'b0000101000110111110 : color = 12'hf00;
15'b0000101000110111111 : color = 12'hf63;
15'b0000101000111000000 : color = 12'he73;
15'b0000101000111000001 : color = 12'he73;
15'b0000101000111000010 : color = 12'he61;
15'b0000101000111000011 : color = 12'hf00;
15'b0000101000111000100 : color = 12'hf53;
15'b0000101000111000101 : color = 12'he73;
15'b0000101000111000110 : color = 12'hf51;
15'b0000101000111000111 : color = 12'hf10;
15'b0000101000111001000 : color = 12'hf52;
15'b0000101000111001001 : color = 12'he72;
15'b0000101000111001010 : color = 12'hf10;
15'b0000101000111001011 : color = 12'hf32;
15'b0000101000111001100 : color = 12'he73;
15'b0000101000111001101 : color = 12'he73;
15'b0000101000111001110 : color = 12'he73;
15'b0000101000111001111 : color = 12'he72;
15'b0000101000111010000 : color = 12'hf10;
15'b0000101000111010001 : color = 12'hf32;
15'b0000101000111010010 : color = 12'he73;
15'b0000101000111010011 : color = 12'he73;
15'b0000101000111010100 : color = 12'he73;
15'b0000101000111010101 : color = 12'he73;
15'b0000101000111010110 : color = 12'he73;
15'b0000101000111010111 : color = 12'he73;
15'b0000101000111011000 : color = 12'he73;
15'b0000101000111011001 : color = 12'he73;
15'b0000101000111011010 : color = 12'he73;
15'b0000101000111011011 : color = 12'he73;
15'b0000101000111011100 : color = 12'he73;
15'b0000101000111011101 : color = 12'he73;
15'b0000101000111011110 : color = 12'he73;
15'b0000101000111011111 : color = 12'he73;
15'b0000101000111100000 : color = 12'he73;
15'b0000101000111100001 : color = 12'he73;
15'b0000101000111100010 : color = 12'he73;
15'b0000101000111100011 : color = 12'he73;
15'b0000101000111100100 : color = 12'he73;
15'b0000101000111100101 : color = 12'he73;
15'b0000101000111100110 : color = 12'he73;
15'b0000101000111100111 : color = 12'he73;
15'b0000101000111101000 : color = 12'he73;
15'b0000101000111101001 : color = 12'he73;
15'b0000101000111101010 : color = 12'he73;
15'b0000101000111101011 : color = 12'he73;
15'b0000101000111101100 : color = 12'he73;
15'b0000101000111101101 : color = 12'he73;
15'b0000101000111101110 : color = 12'he73;
15'b0000101000111101111 : color = 12'hf40;
15'b0000101000111110000 : color = 12'hf00;
15'b0000101000111110001 : color = 12'hf31;
15'b0000101000111110010 : color = 12'hf00;
15'b0000101000111110011 : color = 12'hf53;
15'b0000101000111110100 : color = 12'hf40;
15'b0000101000111110101 : color = 12'hf53;
15'b0000101000111110110 : color = 12'he73;
15'b0000101000111110111 : color = 12'he73;
15'b0000101000111111000 : color = 12'he73;
15'b0000101000111111001 : color = 12'he73;
15'b0000101000111111010 : color = 12'he73;
15'b0000101000111111011 : color = 12'he73;
15'b0000101000111111100 : color = 12'he73;
15'b0000101000111111101 : color = 12'he73;
15'b0000101000111111110 : color = 12'he73;
15'b0000101000111111111 : color = 12'he73;
15'b0000101001000000000 : color = 12'he73;
15'b0000101001000000001 : color = 12'he73;
15'b0000101001000000010 : color = 12'he73;
15'b0000101001000000011 : color = 12'he73;
15'b0000101001000000100 : color = 12'he73;
15'b0000101001000000101 : color = 12'he73;
15'b0000101001000000110 : color = 12'he73;
15'b0000101001000000111 : color = 12'he73;
15'b0000101001000001000 : color = 12'he73;
15'b0000101001000001001 : color = 12'he73;
15'b0000101001000001010 : color = 12'he73;
15'b0000101001000001011 : color = 12'he73;
15'b0000101001000001100 : color = 12'he73;
15'b0000101001000001101 : color = 12'he73;
15'b0000101001000001110 : color = 12'he73;
15'b0000101001000001111 : color = 12'he73;
15'b0000101001000010000 : color = 12'he73;
15'b0000101001000010001 : color = 12'he73;
15'b0000101001000010010 : color = 12'he73;
15'b0000101001000010011 : color = 12'he73;
15'b0000101001000010100 : color = 12'he73;
15'b0000101001000010101 : color = 12'he73;
15'b0000101001000010110 : color = 12'he73;
15'b0000101001000010111 : color = 12'he73;
15'b0000101001000011000 : color = 12'he72;
15'b0000101001000011001 : color = 12'hf00;
15'b0000101001000011010 : color = 12'hf42;
15'b0000101001000011011 : color = 12'he73;
15'b0000101001000011100 : color = 12'he73;
15'b0000101001000011101 : color = 12'he73;
15'b0000101001000011110 : color = 12'hf40;
15'b0000101001000011111 : color = 12'hf42;
15'b0000101001000100000 : color = 12'he73;
15'b0000101001000100001 : color = 12'he73;
15'b0000101001000100010 : color = 12'he72;
15'b0000101001000100011 : color = 12'hf10;
15'b0000101001000100100 : color = 12'hf32;
15'b0000101001000100101 : color = 12'he73;
15'b0000101001000100110 : color = 12'he73;
15'b0000101001000100111 : color = 12'he73;
15'b0000101001000101000 : color = 12'hf40;
15'b0000101001000101001 : color = 12'hf01;
15'b0000101001000101010 : color = 12'hf73;
15'b0000101001000101011 : color = 12'he73;
15'b0000101001000101100 : color = 12'he73;
15'b0000101001000101101 : color = 12'he73;
15'b0000101001000101110 : color = 12'he73;
15'b0000101001000101111 : color = 12'he73;
15'b0000101001000110000 : color = 12'he73;
15'b0000101001000110001 : color = 12'he73;
15'b0000101001000110010 : color = 12'he73;
15'b0000101001000110011 : color = 12'he73;
15'b0000101001000110100 : color = 12'he73;
15'b0000101001000110101 : color = 12'he73;
15'b0000101001000110110 : color = 12'he73;
15'b0000101001000110111 : color = 12'he73;
15'b0000101001000111000 : color = 12'he73;
15'b0000101001000111001 : color = 12'he73;
15'b0000101001000111010 : color = 12'he73;
15'b0000101001000111011 : color = 12'he73;
15'b0000101001000111100 : color = 12'he73;
15'b0000101001000111101 : color = 12'he73;
15'b0000101001000111110 : color = 12'he73;
15'b0000101001000111111 : color = 12'he73;
15'b0000101001001000000 : color = 12'he73;
15'b0000101001001000001 : color = 12'he73;
15'b0000101001001000010 : color = 12'he73;
15'b0000101001001000011 : color = 12'he73;
15'b0000101001001000100 : color = 12'he73;
15'b0000101001001000101 : color = 12'he73;
15'b0000101001001000110 : color = 12'he61;
15'b0000101001001000111 : color = 12'hf32;
15'b0000101001001001000 : color = 12'he73;
15'b0000101001001001001 : color = 12'he73;
15'b0000101001001001010 : color = 12'he73;
15'b0000101001001001011 : color = 12'he73;
15'b0000101001001001100 : color = 12'hf40;
15'b0000101001001001101 : color = 12'hf00;
15'b0000101001001001110 : color = 12'hf53;
15'b0000101001001001111 : color = 12'he73;
15'b0000101001001010000 : color = 12'he73;
15'b0000101001001010001 : color = 12'he73;
15'b0000101001001010010 : color = 12'he73;
15'b0000101001001010011 : color = 12'he73;
15'b0000101001001010100 : color = 12'he73;
15'b0000101001001010101 : color = 12'he73;
15'b0000101001001010110 : color = 12'he73;
15'b0000101001001010111 : color = 12'he73;
15'b0000101001001011000 : color = 12'he73;
15'b0000101001001011001 : color = 12'he73;
15'b0000101001001011010 : color = 12'he73;
15'b0000101001001011011 : color = 12'he73;
15'b0000101001001011100 : color = 12'he73;
15'b0000101001001011101 : color = 12'he73;
15'b0000101001001011110 : color = 12'he73;
15'b0000101001001011111 : color = 12'he73;
15'b0000101001001100000 : color = 12'he73;
15'b0000101001001100001 : color = 12'he73;
15'b0000101001001100010 : color = 12'he73;
15'b0000101001001100011 : color = 12'he73;
15'b0000101001001100100 : color = 12'he73;
15'b0000101001001100101 : color = 12'he73;
15'b0000101001001100110 : color = 12'he73;
15'b0000101001001100111 : color = 12'he73;
15'b0000101001001101000 : color = 12'he73;
15'b0000101001001101001 : color = 12'he73;
15'b0000101001001101010 : color = 12'he73;
15'b0000101001001101011 : color = 12'he73;
15'b0000101001001101100 : color = 12'he73;
15'b0000101001001101101 : color = 12'he51;
15'b0000101001001101110 : color = 12'hf00;
15'b0000101001001101111 : color = 12'hf63;
15'b0000101001001110000 : color = 12'he73;
15'b0000101001001110001 : color = 12'he73;
15'b0000101001001110010 : color = 12'hf40;
15'b0000101001001110011 : color = 12'hf00;
15'b0000101001001110100 : color = 12'hf31;
15'b0000101001001110101 : color = 12'hf31;
15'b0000101001001110110 : color = 12'hf31;
15'b0000101001001110111 : color = 12'hf31;
15'b0000101001001111000 : color = 12'hf30;
15'b0000101001001111001 : color = 12'hf00;
15'b0000101001001111010 : color = 12'hf11;
15'b0000101001001111011 : color = 12'hf31;
15'b0000101001001111100 : color = 12'hf31;
15'b0000101001001111101 : color = 12'hf31;
15'b0000101001001111110 : color = 12'hf31;
15'b0000101001001111111 : color = 12'hf10;
15'b0000101001010000000 : color = 12'hf00;
15'b0000101001010000001 : color = 12'hf63;
15'b0000101001010000010 : color = 12'he73;
15'b0000101001010000011 : color = 12'he73;
15'b0000101001010000100 : color = 12'he73;
15'b0000101001010000101 : color = 12'he73;
15'b0000101001010000110 : color = 12'he73;
15'b0000101001010000111 : color = 12'he73;
15'b0000101001010001000 : color = 12'he73;
15'b0000101001010001001 : color = 12'he73;
15'b0000101001010001010 : color = 12'he73;
15'b0000101001010001011 : color = 12'he73;
15'b0000101001010001100 : color = 12'he73;
15'b0000101001010001101 : color = 12'he73;
15'b0000101001010001110 : color = 12'he73;
15'b0000101001010001111 : color = 12'he73;
15'b0000101001010010000 : color = 12'he73;
15'b0000101001010010001 : color = 12'he73;
15'b0000101001010010010 : color = 12'he73;
15'b0000101001010010011 : color = 12'he73;
15'b0000101001010010100 : color = 12'he73;
15'b0000101001010010101 : color = 12'he73;
15'b0000101001010010110 : color = 12'he73;
15'b0000101001010010111 : color = 12'he73;
15'b0000101001010011000 : color = 12'he73;
15'b0000101001010011001 : color = 12'he73;
15'b0000101001010011010 : color = 12'hf30;
15'b0000101001010011011 : color = 12'hf11;
15'b0000101001010011100 : color = 12'hf73;
15'b0000101001010011101 : color = 12'he73;
15'b0000101001010011110 : color = 12'he73;
15'b0000101001010011111 : color = 12'he73;
15'b0000101001010100000 : color = 12'he73;
15'b0000101001010100001 : color = 12'he73;
15'b0000101001010100010 : color = 12'he73;
15'b0000101001010100011 : color = 12'he73;
15'b0000101001010100100 : color = 12'he73;
15'b0000101001010100101 : color = 12'he73;
15'b0000101001010100110 : color = 12'he51;
15'b0000101001010100111 : color = 12'hf00;
15'b0000101001010101000 : color = 12'hf53;
15'b0000101001010101001 : color = 12'he73;
15'b0000101001010101010 : color = 12'he73;
15'b0000101001010101011 : color = 12'he73;
15'b0000101001010101100 : color = 12'he73;
15'b0000101001010101101 : color = 12'he73;
15'b0000101001010101110 : color = 12'he73;
15'b0000101001010101111 : color = 12'he73;
15'b0000101001010110000 : color = 12'he73;
15'b0000101001010110001 : color = 12'he73;
15'b0000101001010110010 : color = 12'he73;
15'b0000101001010110011 : color = 12'he73;
15'b0000101001010110100 : color = 12'he73;
15'b0000101001010110101 : color = 12'he73;
15'b0000101001010110110 : color = 12'he73;
15'b0000101001010110111 : color = 12'he73;
15'b0000101001010111000 : color = 12'he73;
15'b0000101001010111001 : color = 12'he73;
15'b0000101001010111010 : color = 12'he73;
15'b0000101001010111011 : color = 12'he73;
15'b0000101001010111100 : color = 12'he73;
15'b0000101001010111101 : color = 12'he73;
15'b0000101001010111110 : color = 12'he73;
15'b0000101001010111111 : color = 12'he73;
15'b0000101001011000000 : color = 12'he73;
15'b0000101001011000001 : color = 12'he73;
15'b0000101001011000010 : color = 12'he73;
15'b0000101001011000011 : color = 12'he73;
15'b0000101001011000100 : color = 12'he73;
15'b0000101001011000101 : color = 12'he73;
15'b0000101001011000110 : color = 12'he73;
15'b0000101001011000111 : color = 12'hf30;
15'b0000101001011001000 : color = 12'hf11;
15'b0000101001011001001 : color = 12'hf73;
15'b0000101001011001010 : color = 12'he73;
15'b0000101001011001011 : color = 12'he73;
15'b0000101001011001100 : color = 12'he73;
15'b0000101001011001101 : color = 12'he73;
15'b0000101001011001110 : color = 12'he73;
15'b0000101001011001111 : color = 12'he73;
15'b0000101001011010000 : color = 12'he73;
15'b0000101001011010001 : color = 12'he73;
15'b0000101001011010010 : color = 12'he72;
15'b0000101001011010011 : color = 12'hf10;
15'b0000101001011010100 : color = 12'hf32;
15'b0000101001011010101 : color = 12'he73;
15'b0000101001011010110 : color = 12'he73;
15'b0000101001011010111 : color = 12'he73;
15'b0000101001011011000 : color = 12'he73;
15'b0000101001011011001 : color = 12'he73;
15'b0000101001011011010 : color = 12'he73;
15'b0000101001011011011 : color = 12'he73;
15'b0000101001011011100 : color = 12'he73;
15'b0000101001011011101 : color = 12'he73;
15'b0000101001011011110 : color = 12'he73;
15'b0000101001011011111 : color = 12'he73;
15'b0000101001011100000 : color = 12'he73;
15'b0000101001011100001 : color = 12'he73;
15'b0000101001011100010 : color = 12'he73;
15'b0000101001011100011 : color = 12'he73;
15'b0000101001011100100 : color = 12'he73;
15'b0000101001011100101 : color = 12'he73;
15'b0000101001011100110 : color = 12'he73;
15'b0000101001011100111 : color = 12'he73;
15'b0000101001011101000 : color = 12'he73;
15'b0000101001011101001 : color = 12'he73;
15'b0000101001011101010 : color = 12'he73;
15'b0000101001011101011 : color = 12'he73;
15'b0000101001011101100 : color = 12'he73;
15'b0000101001011101101 : color = 12'he73;
15'b0000101001011101110 : color = 12'he73;
15'b0000101001011101111 : color = 12'he73;
15'b0000101001011110000 : color = 12'he73;
15'b0000101001011110001 : color = 12'he72;
15'b0000101001011110010 : color = 12'hf10;
15'b0000101001011110011 : color = 12'hf32;
15'b0000101001011110100 : color = 12'he73;
15'b0000101001011110101 : color = 12'he73;
15'b0000101001011110110 : color = 12'he73;
15'b0000101001011110111 : color = 12'he73;
15'b0000101001011111000 : color = 12'he62;
15'b0000101001011111001 : color = 12'hf52;
15'b0000101001011111010 : color = 12'he73;
15'b0000101001011111011 : color = 12'he73;
15'b0000101001011111100 : color = 12'he73;
15'b0000101001011111101 : color = 12'he73;
15'b0000101001011111110 : color = 12'hf30;
15'b0000101001011111111 : color = 12'hf32;
15'b0000101001100000000 : color = 12'he73;
15'b0000101001100000001 : color = 12'he73;
15'b0000101001100000010 : color = 12'he73;
15'b0000101001100000011 : color = 12'he72;
15'b0000101001100000100 : color = 12'hf73;
15'b0000101001100000101 : color = 12'he73;
15'b0000101001100000110 : color = 12'he73;
15'b0000101001100000111 : color = 12'he73;
15'b0000101001100001000 : color = 12'he73;
15'b0000101001100001001 : color = 12'he73;
15'b0000101001100001010 : color = 12'he73;
15'b0000101001100001011 : color = 12'he73;
15'b0000101001100001100 : color = 12'he73;
15'b0000101001100001101 : color = 12'he73;
15'b0000101001100001110 : color = 12'he73;
15'b0000101001100001111 : color = 12'he73;
15'b0000101001100010000 : color = 12'he73;
15'b0000101001100010001 : color = 12'he73;
15'b0000101001100010010 : color = 12'he73;
15'b0000101001100010011 : color = 12'he73;
15'b0000101001100010100 : color = 12'he73;
15'b0000101001100010101 : color = 12'he73;
15'b0000101001100010110 : color = 12'he73;
15'b0000101001100010111 : color = 12'he73;
15'b0000101001100011000 : color = 12'he73;
15'b0000101001100011001 : color = 12'he73;
15'b0000101001100011010 : color = 12'he73;
15'b0000101001100011011 : color = 12'he73;
15'b0000101001100011100 : color = 12'he73;
15'b0000101001100011101 : color = 12'hf40;
15'b0000101001100011110 : color = 12'hf00;
15'b0000101001100011111 : color = 12'hf00;
15'b0000101001100100000 : color = 12'hf00;
15'b0000101001100100001 : color = 12'hf31;
15'b0000101001100100010 : color = 12'hf30;
15'b0000101001100100011 : color = 12'hf10;
15'b0000101001100100100 : color = 12'hf10;
15'b0000101001100100101 : color = 12'hf10;
15'b0000101001100100110 : color = 12'hf00;
15'b0000101001100100111 : color = 12'hf00;
15'b0000101001100101000 : color = 12'hf00;
15'b0000101001100101001 : color = 12'hf31;
15'b0000101001100101010 : color = 12'hf31;
15'b0000101001100101011 : color = 12'hf31;
15'b0000101001100101100 : color = 12'hf52;
15'b0000101001100101101 : color = 12'hf52;
15'b0000101001100101110 : color = 12'hf41;
15'b0000101001100101111 : color = 12'hf00;
15'b0000101001100110000 : color = 12'hf00;
15'b0000101001100110001 : color = 12'hf53;
15'b0000101001100110010 : color = 12'he73;
15'b0000101001100110011 : color = 12'he73;
15'b0000101001100110100 : color = 12'he73;
15'b0000101001100110101 : color = 12'he73;
15'b0000101001100110110 : color = 12'he73;
15'b0000101001100110111 : color = 12'he73;
15'b0000101001100111000 : color = 12'he73;
15'b0000101001100111001 : color = 12'he73;
15'b0000101001100111010 : color = 12'he73;
15'b0000101001100111011 : color = 12'he73;
15'b0000101001100111100 : color = 12'he73;
15'b0000101001100111101 : color = 12'he73;
15'b0000101001100111110 : color = 12'he73;
15'b0000101001100111111 : color = 12'he73;
15'b0000101001101000000 : color = 12'he73;
15'b0000101001101000001 : color = 12'he73;
15'b0000101001101000010 : color = 12'he73;
15'b0000101001101000011 : color = 12'he73;
15'b0000101001101000100 : color = 12'he73;
15'b0000101001101000101 : color = 12'he73;
15'b0000101001101000110 : color = 12'he61;
15'b0000101001101000111 : color = 12'hf10;
15'b0000101001101001000 : color = 12'hf11;
15'b0000101001101001001 : color = 12'hf52;
15'b0000101001101001010 : color = 12'hf41;
15'b0000101001101001011 : color = 12'hf31;
15'b0000101001101001100 : color = 12'hf10;
15'b0000101001101001101 : color = 12'hf10;
15'b0000101001101001110 : color = 12'hf31;
15'b0000101001101001111 : color = 12'hf52;
15'b0000101001101010000 : color = 12'hf73;
15'b0000101001101010001 : color = 12'he73;
15'b0000101001101010010 : color = 12'he73;
15'b0000101001101010011 : color = 12'he61;
15'b0000101001101010100 : color = 12'hf00;
15'b0000101001101010101 : color = 12'hf42;
15'b0000101001101010110 : color = 12'he73;
15'b0000101001101010111 : color = 12'he73;
15'b0000101001101011000 : color = 12'hf30;
15'b0000101001101011001 : color = 12'hf11;
15'b0000101001101011010 : color = 12'hf73;
15'b0000101001101011011 : color = 12'he73;
15'b0000101001101011100 : color = 12'he73;
15'b0000101001101011101 : color = 12'he73;
15'b0000101001101011110 : color = 12'he73;
15'b0000101001101011111 : color = 12'he73;
15'b0000101001101100000 : color = 12'he73;
15'b0000101001101100001 : color = 12'he73;
15'b0000101001101100010 : color = 12'he73;
15'b0000101001101100011 : color = 12'he73;
15'b0000101001101100100 : color = 12'he73;
15'b0000101001101100101 : color = 12'he73;
15'b0000101001101100110 : color = 12'he73;
15'b0000101001101100111 : color = 12'he73;
15'b0000101001101101000 : color = 12'he73;
15'b0000101001101101001 : color = 12'he73;
15'b0000101001101101010 : color = 12'he73;
15'b0000101001101101011 : color = 12'he73;
15'b0000101001101101100 : color = 12'he73;
15'b0000101001101101101 : color = 12'he73;
15'b0000101001101101110 : color = 12'he73;
15'b0000101001101101111 : color = 12'he73;
15'b0000101000110101110 : color = 12'he73;
15'b0000101000110101111 : color = 12'he73;
15'b0000101000110110000 : color = 12'he73;
15'b0000101000110110001 : color = 12'he73;
15'b0000101000110110010 : color = 12'he73;
15'b0000101000110110011 : color = 12'he73;
15'b0000101000110110100 : color = 12'he73;
15'b0000101000110110101 : color = 12'he73;
15'b0000101000110110110 : color = 12'he73;
15'b0000101000110110111 : color = 12'he73;
15'b0000101000110111000 : color = 12'he73;
15'b0000101000110111001 : color = 12'he73;
15'b0000101000110111010 : color = 12'he72;
15'b0000101000110111011 : color = 12'hf00;
15'b0000101000110111100 : color = 12'hf42;
15'b0000101000110111101 : color = 12'he51;
15'b0000101000110111110 : color = 12'hf00;
15'b0000101000110111111 : color = 12'hf11;
15'b0000101000111000000 : color = 12'hf73;
15'b0000101000111000001 : color = 12'he73;
15'b0000101000111000010 : color = 12'he73;
15'b0000101000111000011 : color = 12'he73;
15'b0000101000111000100 : color = 12'he73;
15'b0000101000111000101 : color = 12'he61;
15'b0000101000111000110 : color = 12'hf00;
15'b0000101000111000111 : color = 12'hf53;
15'b0000101000111001000 : color = 12'he73;
15'b0000101000111001001 : color = 12'hf30;
15'b0000101000111001010 : color = 12'hf53;
15'b0000101000111001011 : color = 12'he73;
15'b0000101000111001100 : color = 12'he73;
15'b0000101000111001101 : color = 12'he73;
15'b0000101000111001110 : color = 12'he73;
15'b0000101000111001111 : color = 12'he73;
15'b0000101000111010000 : color = 12'he73;
15'b0000101000111010001 : color = 12'he73;
15'b0000101000111010010 : color = 12'he73;
15'b0000101000111010011 : color = 12'he73;
15'b0000101000111010100 : color = 12'he73;
15'b0000101000111010101 : color = 12'he73;
15'b0000101000111010110 : color = 12'he73;
15'b0000101000111010111 : color = 12'he73;
15'b0000101000111011000 : color = 12'he73;
15'b0000101000111011001 : color = 12'he73;
15'b0000101000111011010 : color = 12'he73;
15'b0000101000111011011 : color = 12'he73;
15'b0000101000111011100 : color = 12'he73;
15'b0000101000111011101 : color = 12'he73;
15'b0000101000111011110 : color = 12'he73;
15'b0000101000111011111 : color = 12'he73;
15'b0000101000111100000 : color = 12'he73;
15'b0000101000111100001 : color = 12'he73;
15'b0000101000111100010 : color = 12'he73;
15'b0000101000111100011 : color = 12'he73;
15'b0000101000111100100 : color = 12'he73;
15'b0000101000111100101 : color = 12'he73;
15'b0000101000111100110 : color = 12'he51;
15'b0000101000111100111 : color = 12'hf00;
15'b0000101000111101000 : color = 12'hf63;
15'b0000101000111101001 : color = 12'he73;
15'b0000101000111101010 : color = 12'he73;
15'b0000101000111101011 : color = 12'he61;
15'b0000101000111101100 : color = 12'hf00;
15'b0000101000111101101 : color = 12'hf31;
15'b0000101000111101110 : color = 12'hf00;
15'b0000101000111101111 : color = 12'hf11;
15'b0000101000111110000 : color = 12'hf63;
15'b0000101000111110001 : color = 12'he73;
15'b0000101000111110010 : color = 12'he72;
15'b0000101000111110011 : color = 12'hf10;
15'b0000101000111110100 : color = 12'hf32;
15'b0000101000111110101 : color = 12'he73;
15'b0000101000111110110 : color = 12'he73;
15'b0000101000111110111 : color = 12'he73;
15'b0000101000111111000 : color = 12'he72;
15'b0000101000111111001 : color = 12'hf10;
15'b0000101000111111010 : color = 12'hf32;
15'b0000101000111111011 : color = 12'he73;
15'b0000101000111111100 : color = 12'he73;
15'b0000101000111111101 : color = 12'he73;
15'b0000101000111111110 : color = 12'he73;
15'b0000101000111111111 : color = 12'he73;
15'b0000101001000000000 : color = 12'he73;
15'b0000101001000000001 : color = 12'he73;
15'b0000101001000000010 : color = 12'he73;
15'b0000101001000000011 : color = 12'he73;
15'b0000101001000000100 : color = 12'he73;
15'b0000101001000000101 : color = 12'he73;
15'b0000101001000000110 : color = 12'he73;
15'b0000101001000000111 : color = 12'he73;
15'b0000101001000001000 : color = 12'he73;
15'b0000101001000001001 : color = 12'he73;
15'b0000101001000001010 : color = 12'he73;
15'b0000101001000001011 : color = 12'he73;
15'b0000101001000001100 : color = 12'he73;
15'b0000101001000001101 : color = 12'he73;
15'b0000101001000001110 : color = 12'he73;
15'b0000101001000001111 : color = 12'he73;
15'b0000101001000010000 : color = 12'he73;
15'b0000101001000010001 : color = 12'he73;
15'b0000101001000010010 : color = 12'he73;
15'b0000101001000010011 : color = 12'he73;
15'b0000101001000010100 : color = 12'he73;
15'b0000101001000010101 : color = 12'he73;
15'b0000101001000010110 : color = 12'he73;
15'b0000101001000010111 : color = 12'he61;
15'b0000101001000011000 : color = 12'hf00;
15'b0000101001000011001 : color = 12'hf32;
15'b0000101001000011010 : color = 12'he51;
15'b0000101001000011011 : color = 12'hf00;
15'b0000101001000011100 : color = 12'hf53;
15'b0000101001000011101 : color = 12'he72;
15'b0000101001000011110 : color = 12'hf11;
15'b0000101001000011111 : color = 12'hf73;
15'b0000101001000100000 : color = 12'he73;
15'b0000101001000100001 : color = 12'he73;
15'b0000101001000100010 : color = 12'he73;
15'b0000101001000100011 : color = 12'he73;
15'b0000101001000100100 : color = 12'he73;
15'b0000101001000100101 : color = 12'he73;
15'b0000101001000100110 : color = 12'he73;
15'b0000101001000100111 : color = 12'he73;
15'b0000101001000101000 : color = 12'he73;
15'b0000101001000101001 : color = 12'he73;
15'b0000101001000101010 : color = 12'he73;
15'b0000101001000101011 : color = 12'he73;
15'b0000101001000101100 : color = 12'he73;
15'b0000101001000101101 : color = 12'he73;
15'b0000101001000101110 : color = 12'he73;
15'b0000101001000101111 : color = 12'he73;
15'b0000101001000110000 : color = 12'he73;
15'b0000101001000110001 : color = 12'he73;
15'b0000101001000110010 : color = 12'he73;
15'b0000101001000110011 : color = 12'he73;
15'b0000101001000110100 : color = 12'he73;
15'b0000101001000110101 : color = 12'he73;
15'b0000101001000110110 : color = 12'he73;
15'b0000101001000110111 : color = 12'he73;
15'b0000101001000111000 : color = 12'he73;
15'b0000101001000111001 : color = 12'he73;
15'b0000101001000111010 : color = 12'he73;
15'b0000101001000111011 : color = 12'he61;
15'b0000101001000111100 : color = 12'hf31;
15'b0000101001000111101 : color = 12'hf31;
15'b0000101001000111110 : color = 12'hf31;
15'b0000101001000111111 : color = 12'hf31;
15'b0000101001001000000 : color = 12'hf31;
15'b0000101001001000001 : color = 12'hf30;
15'b0000101001001000010 : color = 12'hf00;
15'b0000101001001000011 : color = 12'hf11;
15'b0000101001001000100 : color = 12'hf31;
15'b0000101001001000101 : color = 12'hf31;
15'b0000101001001000110 : color = 12'hf30;
15'b0000101001001000111 : color = 12'hf00;
15'b0000101001001001000 : color = 12'hf00;
15'b0000101001001001001 : color = 12'hf42;
15'b0000101001001001010 : color = 12'he73;
15'b0000101001001001011 : color = 12'he72;
15'b0000101001001001100 : color = 12'hf10;
15'b0000101001001001101 : color = 12'hf32;
15'b0000101001001001110 : color = 12'he73;
15'b0000101001001001111 : color = 12'he73;
15'b0000101001001010000 : color = 12'he73;
15'b0000101001001010001 : color = 12'hf40;
15'b0000101001001010010 : color = 12'hf01;
15'b0000101001001010011 : color = 12'hf73;
15'b0000101001001010100 : color = 12'he73;
15'b0000101001001010101 : color = 12'he73;
15'b0000101001001010110 : color = 12'he73;
15'b0000101001001010111 : color = 12'he73;
15'b0000101001001011000 : color = 12'he73;
15'b0000101001001011001 : color = 12'he73;
15'b0000101001001011010 : color = 12'he73;
15'b0000101001001011011 : color = 12'he73;
15'b0000101001001011100 : color = 12'he73;
15'b0000101001001011101 : color = 12'he73;
15'b0000101001001011110 : color = 12'he73;
15'b0000101001001011111 : color = 12'he73;
15'b0000101001001100000 : color = 12'he73;
15'b0000101001001100001 : color = 12'he73;
15'b0000101001001100010 : color = 12'he73;
15'b0000101001001100011 : color = 12'he73;
15'b0000101001001100100 : color = 12'he73;
15'b0000101001001100101 : color = 12'he73;
15'b0000101001001100110 : color = 12'he73;
15'b0000101001001100111 : color = 12'he73;
15'b0000101001001101000 : color = 12'he73;
15'b0000101001001101001 : color = 12'he73;
15'b0000101001001101010 : color = 12'he73;
15'b0000101001001101011 : color = 12'he73;
15'b0000101001001101100 : color = 12'he73;
15'b0000101001001101101 : color = 12'he73;
15'b0000101001001101110 : color = 12'he73;
15'b0000101001001101111 : color = 12'he72;
15'b0000101001001110000 : color = 12'hf10;
15'b0000101001001110001 : color = 12'hf53;
15'b0000101001001110010 : color = 12'he73;
15'b0000101001001110011 : color = 12'he73;
15'b0000101001001110100 : color = 12'he72;
15'b0000101001001110101 : color = 12'hf00;
15'b0000101001001110110 : color = 12'hf11;
15'b0000101001001110111 : color = 12'hf73;
15'b0000101001001111000 : color = 12'he73;
15'b0000101001001111001 : color = 12'he73;
15'b0000101001001111010 : color = 12'he73;
15'b0000101001001111011 : color = 12'he73;
15'b0000101001001111100 : color = 12'he73;
15'b0000101001001111101 : color = 12'he73;
15'b0000101001001111110 : color = 12'he73;
15'b0000101001001111111 : color = 12'he73;
15'b0000101001010000000 : color = 12'he73;
15'b0000101001010000001 : color = 12'he73;
15'b0000101001010000010 : color = 12'he73;
15'b0000101001010000011 : color = 12'he73;
15'b0000101001010000100 : color = 12'he73;
15'b0000101001010000101 : color = 12'he73;
15'b0000101001010000110 : color = 12'he73;
15'b0000101001010000111 : color = 12'he73;
15'b0000101001010001000 : color = 12'he73;
15'b0000101001010001001 : color = 12'he73;
15'b0000101001010001010 : color = 12'he73;
15'b0000101001010001011 : color = 12'he73;
15'b0000101001010001100 : color = 12'he73;
15'b0000101001010001101 : color = 12'he73;
15'b0000101001010001110 : color = 12'he73;
15'b0000101001010001111 : color = 12'he73;
15'b0000101001010010000 : color = 12'he73;
15'b0000101001010010001 : color = 12'he73;
15'b0000101001010010010 : color = 12'he73;
15'b0000101001010010011 : color = 12'he73;
15'b0000101001010010100 : color = 12'he73;
15'b0000101001010010101 : color = 12'he73;
15'b0000101001010010110 : color = 12'he51;
15'b0000101001010010111 : color = 12'hf00;
15'b0000101001010011000 : color = 12'hf63;
15'b0000101001010011001 : color = 12'he73;
15'b0000101001010011010 : color = 12'he73;
15'b0000101001010011011 : color = 12'hf30;
15'b0000101001010011100 : color = 12'hf11;
15'b0000101001010011101 : color = 12'hf73;
15'b0000101001010011110 : color = 12'he73;
15'b0000101001010011111 : color = 12'he73;
15'b0000101001010100000 : color = 12'he73;
15'b0000101001010100001 : color = 12'he61;
15'b0000101001010100010 : color = 12'hf00;
15'b0000101001010100011 : color = 12'hf53;
15'b0000101001010100100 : color = 12'he73;
15'b0000101001010100101 : color = 12'he73;
15'b0000101001010100110 : color = 12'he73;
15'b0000101001010100111 : color = 12'he73;
15'b0000101001010101000 : color = 12'he51;
15'b0000101001010101001 : color = 12'hf00;
15'b0000101001010101010 : color = 12'hf63;
15'b0000101001010101011 : color = 12'he73;
15'b0000101001010101100 : color = 12'he73;
15'b0000101001010101101 : color = 12'he73;
15'b0000101001010101110 : color = 12'he73;
15'b0000101001010101111 : color = 12'he73;
15'b0000101001010110000 : color = 12'he73;
15'b0000101001010110001 : color = 12'he73;
15'b0000101001010110010 : color = 12'he73;
15'b0000101001010110011 : color = 12'he73;
15'b0000101001010110100 : color = 12'he73;
15'b0000101001010110101 : color = 12'he73;
15'b0000101001010110110 : color = 12'he73;
15'b0000101001010110111 : color = 12'he73;
15'b0000101001010111000 : color = 12'he73;
15'b0000101001010111001 : color = 12'he73;
15'b0000101001010111010 : color = 12'he73;
15'b0000101001010111011 : color = 12'he73;
15'b0000101001010111100 : color = 12'he73;
15'b0000101001010111101 : color = 12'he73;
15'b0000101001010111110 : color = 12'he73;
15'b0000101001010111111 : color = 12'he73;
15'b0000101001011000000 : color = 12'he73;
15'b0000101001011000001 : color = 12'he73;
15'b0000101001011000010 : color = 12'he72;
15'b0000101001011000011 : color = 12'hf10;
15'b0000101001011000100 : color = 12'hf32;
15'b0000101001011000101 : color = 12'he73;
15'b0000101001011000110 : color = 12'he73;
15'b0000101001011000111 : color = 12'he73;
15'b0000101001011001000 : color = 12'he73;
15'b0000101001011001001 : color = 12'he73;
15'b0000101001011001010 : color = 12'he73;
15'b0000101001011001011 : color = 12'he73;
15'b0000101001011001100 : color = 12'he73;
15'b0000101001011001101 : color = 12'he73;
15'b0000101001011001110 : color = 12'he73;
15'b0000101001011001111 : color = 12'he51;
15'b0000101001011010000 : color = 12'hf00;
15'b0000101001011010001 : color = 12'hf53;
15'b0000101001011010010 : color = 12'he73;
15'b0000101001011010011 : color = 12'he73;
15'b0000101001011010100 : color = 12'he73;
15'b0000101001011010101 : color = 12'he73;
15'b0000101001011010110 : color = 12'he73;
15'b0000101001011010111 : color = 12'he73;
15'b0000101001011011000 : color = 12'he73;
15'b0000101001011011001 : color = 12'he73;
15'b0000101001011011010 : color = 12'he73;
15'b0000101001011011011 : color = 12'he73;
15'b0000101001011011100 : color = 12'he73;
15'b0000101001011011101 : color = 12'he73;
15'b0000101001011011110 : color = 12'he73;
15'b0000101001011011111 : color = 12'he73;
15'b0000101001011100000 : color = 12'he73;
15'b0000101001011100001 : color = 12'he73;
15'b0000101001011100010 : color = 12'he73;
15'b0000101001011100011 : color = 12'he73;
15'b0000101001011100100 : color = 12'he73;
15'b0000101001011100101 : color = 12'he73;
15'b0000101001011100110 : color = 12'he73;
15'b0000101001011100111 : color = 12'he73;
15'b0000101001011101000 : color = 12'he73;
15'b0000101001011101001 : color = 12'he73;
15'b0000101001011101010 : color = 12'he73;
15'b0000101001011101011 : color = 12'he73;
15'b0000101001011101100 : color = 12'he73;
15'b0000101001011101101 : color = 12'he73;
15'b0000101001011101110 : color = 12'he73;
15'b0000101001011101111 : color = 12'he73;
15'b0000101001011110000 : color = 12'hf30;
15'b0000101001011110001 : color = 12'hf00;
15'b0000101001011110010 : color = 12'hf31;
15'b0000101001011110011 : color = 12'hf31;
15'b0000101001011110100 : color = 12'hf31;
15'b0000101001011110101 : color = 12'hf31;
15'b0000101001011110110 : color = 12'hf31;
15'b0000101001011110111 : color = 12'hf31;
15'b0000101001011111000 : color = 12'hf31;
15'b0000101001011111001 : color = 12'hf31;
15'b0000101001011111010 : color = 12'hf31;
15'b0000101001011111011 : color = 12'hf31;
15'b0000101001011111100 : color = 12'hf00;
15'b0000101001011111101 : color = 12'hf32;
15'b0000101001011111110 : color = 12'he73;
15'b0000101001011111111 : color = 12'he73;
15'b0000101001100000000 : color = 12'he73;
15'b0000101001100000001 : color = 12'he73;
15'b0000101001100000010 : color = 12'he73;
15'b0000101001100000011 : color = 12'he73;
15'b0000101001100000100 : color = 12'he73;
15'b0000101001100000101 : color = 12'he73;
15'b0000101001100000110 : color = 12'he73;
15'b0000101001100000111 : color = 12'he73;
15'b0000101001100001000 : color = 12'he73;
15'b0000101001100001001 : color = 12'he73;
15'b0000101001100001010 : color = 12'he73;
15'b0000101001100001011 : color = 12'he73;
15'b0000101001100001100 : color = 12'he73;
15'b0000101001100001101 : color = 12'he73;
15'b0000101001100001110 : color = 12'he73;
15'b0000101001100001111 : color = 12'he73;
15'b0000101001100010000 : color = 12'he73;
15'b0000101001100010001 : color = 12'he73;
15'b0000101001100010010 : color = 12'he73;
15'b0000101001100010011 : color = 12'he73;
15'b0000101001100010100 : color = 12'he73;
15'b0000101001100010101 : color = 12'he73;
15'b0000101001100010110 : color = 12'he73;
15'b0000101001100010111 : color = 12'he73;
15'b0000101001100011000 : color = 12'he73;
15'b0000101001100011001 : color = 12'he73;
15'b0000101001100011010 : color = 12'he72;
15'b0000101001100011011 : color = 12'hf10;
15'b0000101001100011100 : color = 12'hf32;
15'b0000101001100011101 : color = 12'he73;
15'b0000101001100011110 : color = 12'he73;
15'b0000101001100011111 : color = 12'he73;
15'b0000101001100100000 : color = 12'he73;
15'b0000101001100100001 : color = 12'he73;
15'b0000101001100100010 : color = 12'he73;
15'b0000101001100100011 : color = 12'he73;
15'b0000101001100100100 : color = 12'he73;
15'b0000101001100100101 : color = 12'he73;
15'b0000101001100100110 : color = 12'he73;
15'b0000101001100100111 : color = 12'hf30;
15'b0000101001100101000 : color = 12'hf32;
15'b0000101001100101001 : color = 12'he73;
15'b0000101001100101010 : color = 12'he73;
15'b0000101001100101011 : color = 12'he73;
15'b0000101001100101100 : color = 12'he73;
15'b0000101001100101101 : color = 12'he73;
15'b0000101001100101110 : color = 12'he73;
15'b0000101001100101111 : color = 12'he73;
15'b0000101001100110000 : color = 12'he73;
15'b0000101001100110001 : color = 12'he73;
15'b0000101001100110010 : color = 12'he73;
15'b0000101001100110011 : color = 12'he73;
15'b0000101001100110100 : color = 12'he73;
15'b0000101001100110101 : color = 12'he73;
15'b0000101001100110110 : color = 12'he73;
15'b0000101001100110111 : color = 12'he73;
15'b0000101001100111000 : color = 12'he73;
15'b0000101001100111001 : color = 12'he73;
15'b0000101001100111010 : color = 12'he73;
15'b0000101001100111011 : color = 12'he73;
15'b0000101001100111100 : color = 12'he73;
15'b0000101001100111101 : color = 12'he73;
15'b0000101001100111110 : color = 12'he73;
15'b0000101001100111111 : color = 12'he73;
15'b0000101001101000000 : color = 12'he73;
15'b0000101001101000001 : color = 12'he73;
15'b0000101001101000010 : color = 12'he73;
15'b0000101001101000011 : color = 12'he73;
15'b0000101001101000100 : color = 12'he73;
15'b0000101001101000101 : color = 12'he73;
15'b0000101001101000110 : color = 12'he72;
15'b0000101001101000111 : color = 12'hf00;
15'b0000101001101001000 : color = 12'hf00;
15'b0000101001101001001 : color = 12'hf00;
15'b0000101001101001010 : color = 12'hf31;
15'b0000101001101001011 : color = 12'hf52;
15'b0000101001101001100 : color = 12'hf62;
15'b0000101001101001101 : color = 12'hf62;
15'b0000101001101001110 : color = 12'he73;
15'b0000101001101001111 : color = 12'he51;
15'b0000101001101010000 : color = 12'hf00;
15'b0000101001101010001 : color = 12'hf53;
15'b0000101001101010010 : color = 12'he73;
15'b0000101001101010011 : color = 12'he73;
15'b0000101001101010100 : color = 12'he73;
15'b0000101001101010101 : color = 12'he73;
15'b0000101001101010110 : color = 12'he73;
15'b0000101001101010111 : color = 12'he73;
15'b0000101001101011000 : color = 12'hf40;
15'b0000101001101011001 : color = 12'hf00;
15'b0000101001101011010 : color = 12'hf53;
15'b0000101001101011011 : color = 12'he73;
15'b0000101001101011100 : color = 12'he73;
15'b0000101001101011101 : color = 12'he73;
15'b0000101001101011110 : color = 12'he73;
15'b0000101001101011111 : color = 12'he73;
15'b0000101001101100000 : color = 12'he73;
15'b0000101001101100001 : color = 12'he73;
15'b0000101001101100010 : color = 12'he73;
15'b0000101001101100011 : color = 12'he73;
15'b0000101001101100100 : color = 12'he73;
15'b0000101001101100101 : color = 12'he73;
15'b0000101001101100110 : color = 12'he73;
15'b0000101001101100111 : color = 12'he73;
15'b0000101001101101000 : color = 12'he73;
15'b0000101001101101001 : color = 12'he73;
15'b0000101001101101010 : color = 12'he73;
15'b0000101001101101011 : color = 12'he73;
15'b0000101001101101100 : color = 12'he73;
15'b0000101001101101101 : color = 12'he73;
15'b0000101001101101110 : color = 12'he73;
15'b0000101001101101111 : color = 12'he51;
15'b0000101001101110000 : color = 12'hf00;
15'b0000101001101110001 : color = 12'hf00;
15'b0000101001101110010 : color = 12'hf00;
15'b0000101001101110011 : color = 12'hf11;
15'b0000101001101110100 : color = 12'hf42;
15'b0000101001101110101 : color = 12'hf73;
15'b0000101001101110110 : color = 12'he73;
15'b0000101001101110111 : color = 12'he73;
15'b0000101001101111000 : color = 12'he73;
15'b0000101001101111001 : color = 12'he73;
15'b0000101001101111010 : color = 12'he73;
15'b0000101001101111011 : color = 12'he73;
15'b0000101001101111100 : color = 12'he61;
15'b0000101001101111101 : color = 12'hf00;
15'b0000101001101111110 : color = 12'hf42;
15'b0000101001101111111 : color = 12'he73;
15'b0000101001110000000 : color = 12'he73;
15'b0000101001110000001 : color = 12'hf30;
15'b0000101001110000010 : color = 12'hf11;
15'b0000101001110000011 : color = 12'hf73;
15'b0000101001110000100 : color = 12'he73;
15'b0000101001110000101 : color = 12'he73;
15'b0000101001110000110 : color = 12'he73;
15'b0000101001110000111 : color = 12'he73;
15'b0000101001110001000 : color = 12'he73;
15'b0000101001110001001 : color = 12'he73;
15'b0000101001110001010 : color = 12'he73;
15'b0000101001110001011 : color = 12'he73;
15'b0000101001110001100 : color = 12'he73;
15'b0000101001110001101 : color = 12'he73;
15'b0000101001110001110 : color = 12'he73;
15'b0000101001110001111 : color = 12'he73;
15'b0000101001110010000 : color = 12'he73;
15'b0000101001110010001 : color = 12'he73;
15'b0000101001110010010 : color = 12'he73;
15'b0000101001110010011 : color = 12'he73;
15'b0000101001110010100 : color = 12'he73;
15'b0000101001110010101 : color = 12'he73;
15'b0000101001110010110 : color = 12'he73;
15'b0000101001110010111 : color = 12'he73;
15'b0000101001110011000 : color = 12'he73;
15'b0000101000111010111 : color = 12'he73;
15'b0000101000111011000 : color = 12'he73;
15'b0000101000111011001 : color = 12'he73;
15'b0000101000111011010 : color = 12'he73;
15'b0000101000111011011 : color = 12'he73;
15'b0000101000111011100 : color = 12'he73;
15'b0000101000111011101 : color = 12'he73;
15'b0000101000111011110 : color = 12'he73;
15'b0000101000111011111 : color = 12'he73;
15'b0000101000111100000 : color = 12'he73;
15'b0000101000111100001 : color = 12'he73;
15'b0000101000111100010 : color = 12'he73;
15'b0000101000111100011 : color = 12'hf40;
15'b0000101000111100100 : color = 12'hf11;
15'b0000101000111100101 : color = 12'hf73;
15'b0000101000111100110 : color = 12'he72;
15'b0000101000111100111 : color = 12'hf10;
15'b0000101000111101000 : color = 12'hf00;
15'b0000101000111101001 : color = 12'hf42;
15'b0000101000111101010 : color = 12'he73;
15'b0000101000111101011 : color = 12'he73;
15'b0000101000111101100 : color = 12'he73;
15'b0000101000111101101 : color = 12'he73;
15'b0000101000111101110 : color = 12'hf40;
15'b0000101000111101111 : color = 12'hf01;
15'b0000101000111110000 : color = 12'hf73;
15'b0000101000111110001 : color = 12'he73;
15'b0000101000111110010 : color = 12'hf40;
15'b0000101000111110011 : color = 12'hf32;
15'b0000101000111110100 : color = 12'he73;
15'b0000101000111110101 : color = 12'he73;
15'b0000101000111110110 : color = 12'he73;
15'b0000101000111110111 : color = 12'he73;
15'b0000101000111111000 : color = 12'he73;
15'b0000101000111111001 : color = 12'he73;
15'b0000101000111111010 : color = 12'he73;
15'b0000101000111111011 : color = 12'he73;
15'b0000101000111111100 : color = 12'he73;
15'b0000101000111111101 : color = 12'he73;
15'b0000101000111111110 : color = 12'he73;
15'b0000101000111111111 : color = 12'he73;
15'b0000101001000000000 : color = 12'he73;
15'b0000101001000000001 : color = 12'he73;
15'b0000101001000000010 : color = 12'he73;
15'b0000101001000000011 : color = 12'he73;
15'b0000101001000000100 : color = 12'he73;
15'b0000101001000000101 : color = 12'he73;
15'b0000101001000000110 : color = 12'he73;
15'b0000101001000000111 : color = 12'he73;
15'b0000101001000001000 : color = 12'he73;
15'b0000101001000001001 : color = 12'he73;
15'b0000101001000001010 : color = 12'he73;
15'b0000101001000001011 : color = 12'he73;
15'b0000101001000001100 : color = 12'he73;
15'b0000101001000001101 : color = 12'he73;
15'b0000101001000001110 : color = 12'he73;
15'b0000101001000001111 : color = 12'he51;
15'b0000101001000010000 : color = 12'hf00;
15'b0000101001000010001 : color = 12'hf63;
15'b0000101001000010010 : color = 12'he73;
15'b0000101001000010011 : color = 12'he73;
15'b0000101001000010100 : color = 12'hf40;
15'b0000101001000010101 : color = 12'hf00;
15'b0000101001000010110 : color = 12'hf00;
15'b0000101001000010111 : color = 12'hf32;
15'b0000101001000011000 : color = 12'he73;
15'b0000101001000011001 : color = 12'he73;
15'b0000101001000011010 : color = 12'he73;
15'b0000101001000011011 : color = 12'he72;
15'b0000101001000011100 : color = 12'hf10;
15'b0000101001000011101 : color = 12'hf32;
15'b0000101001000011110 : color = 12'he62;
15'b0000101001000011111 : color = 12'hf10;
15'b0000101001000100000 : color = 12'hf10;
15'b0000101001000100001 : color = 12'hf10;
15'b0000101001000100010 : color = 12'hf00;
15'b0000101001000100011 : color = 12'hf32;
15'b0000101001000100100 : color = 12'he73;
15'b0000101001000100101 : color = 12'he73;
15'b0000101001000100110 : color = 12'he73;
15'b0000101001000100111 : color = 12'he73;
15'b0000101001000101000 : color = 12'he73;
15'b0000101001000101001 : color = 12'he73;
15'b0000101001000101010 : color = 12'he73;
15'b0000101001000101011 : color = 12'he73;
15'b0000101001000101100 : color = 12'he73;
15'b0000101001000101101 : color = 12'he73;
15'b0000101001000101110 : color = 12'he73;
15'b0000101001000101111 : color = 12'he73;
15'b0000101001000110000 : color = 12'he73;
15'b0000101001000110001 : color = 12'he73;
15'b0000101001000110010 : color = 12'he73;
15'b0000101001000110011 : color = 12'he73;
15'b0000101001000110100 : color = 12'he73;
15'b0000101001000110101 : color = 12'he73;
15'b0000101001000110110 : color = 12'he73;
15'b0000101001000110111 : color = 12'he73;
15'b0000101001000111000 : color = 12'he73;
15'b0000101001000111001 : color = 12'he73;
15'b0000101001000111010 : color = 12'he73;
15'b0000101001000111011 : color = 12'he73;
15'b0000101001000111100 : color = 12'he73;
15'b0000101001000111101 : color = 12'he73;
15'b0000101001000111110 : color = 12'he73;
15'b0000101001000111111 : color = 12'he72;
15'b0000101001001000000 : color = 12'hf10;
15'b0000101001001000001 : color = 12'hf01;
15'b0000101001001000010 : color = 12'hf73;
15'b0000101001001000011 : color = 12'he51;
15'b0000101001001000100 : color = 12'hf00;
15'b0000101001001000101 : color = 12'hf53;
15'b0000101001001000110 : color = 12'he73;
15'b0000101001001000111 : color = 12'hf40;
15'b0000101001001001000 : color = 12'hf11;
15'b0000101001001001001 : color = 12'hf73;
15'b0000101001001001010 : color = 12'he73;
15'b0000101001001001011 : color = 12'he73;
15'b0000101001001001100 : color = 12'he73;
15'b0000101001001001101 : color = 12'he73;
15'b0000101001001001110 : color = 12'he73;
15'b0000101001001001111 : color = 12'he73;
15'b0000101001001010000 : color = 12'he73;
15'b0000101001001010001 : color = 12'he73;
15'b0000101001001010010 : color = 12'he73;
15'b0000101001001010011 : color = 12'he73;
15'b0000101001001010100 : color = 12'he73;
15'b0000101001001010101 : color = 12'he73;
15'b0000101001001010110 : color = 12'he73;
15'b0000101001001010111 : color = 12'he73;
15'b0000101001001011000 : color = 12'he73;
15'b0000101001001011001 : color = 12'he73;
15'b0000101001001011010 : color = 12'he73;
15'b0000101001001011011 : color = 12'he73;
15'b0000101001001011100 : color = 12'he73;
15'b0000101001001011101 : color = 12'he73;
15'b0000101001001011110 : color = 12'he73;
15'b0000101001001011111 : color = 12'he73;
15'b0000101001001100000 : color = 12'he73;
15'b0000101001001100001 : color = 12'he73;
15'b0000101001001100010 : color = 12'he73;
15'b0000101001001100011 : color = 12'he73;
15'b0000101001001100100 : color = 12'he73;
15'b0000101001001100101 : color = 12'he73;
15'b0000101001001100110 : color = 12'he73;
15'b0000101001001100111 : color = 12'he73;
15'b0000101001001101000 : color = 12'he73;
15'b0000101001001101001 : color = 12'he73;
15'b0000101001001101010 : color = 12'he72;
15'b0000101001001101011 : color = 12'hf00;
15'b0000101001001101100 : color = 12'hf42;
15'b0000101001001101101 : color = 12'he73;
15'b0000101001001101110 : color = 12'he73;
15'b0000101001001101111 : color = 12'he73;
15'b0000101001001110000 : color = 12'he73;
15'b0000101001001110001 : color = 12'he73;
15'b0000101001001110010 : color = 12'he73;
15'b0000101001001110011 : color = 12'he73;
15'b0000101001001110100 : color = 12'he72;
15'b0000101001001110101 : color = 12'hf10;
15'b0000101001001110110 : color = 12'hf32;
15'b0000101001001110111 : color = 12'he73;
15'b0000101001001111000 : color = 12'he73;
15'b0000101001001111001 : color = 12'he73;
15'b0000101001001111010 : color = 12'hf40;
15'b0000101001001111011 : color = 12'hf01;
15'b0000101001001111100 : color = 12'hf73;
15'b0000101001001111101 : color = 12'he73;
15'b0000101001001111110 : color = 12'he73;
15'b0000101001001111111 : color = 12'he73;
15'b0000101001010000000 : color = 12'he73;
15'b0000101001010000001 : color = 12'he73;
15'b0000101001010000010 : color = 12'he73;
15'b0000101001010000011 : color = 12'he73;
15'b0000101001010000100 : color = 12'he73;
15'b0000101001010000101 : color = 12'he73;
15'b0000101001010000110 : color = 12'he73;
15'b0000101001010000111 : color = 12'he73;
15'b0000101001010001000 : color = 12'he73;
15'b0000101001010001001 : color = 12'he73;
15'b0000101001010001010 : color = 12'he73;
15'b0000101001010001011 : color = 12'he73;
15'b0000101001010001100 : color = 12'he73;
15'b0000101001010001101 : color = 12'he73;
15'b0000101001010001110 : color = 12'he73;
15'b0000101001010001111 : color = 12'he73;
15'b0000101001010010000 : color = 12'he73;
15'b0000101001010010001 : color = 12'he73;
15'b0000101001010010010 : color = 12'he73;
15'b0000101001010010011 : color = 12'he73;
15'b0000101001010010100 : color = 12'he73;
15'b0000101001010010101 : color = 12'he73;
15'b0000101001010010110 : color = 12'he73;
15'b0000101001010010111 : color = 12'he73;
15'b0000101001010011000 : color = 12'he73;
15'b0000101001010011001 : color = 12'he51;
15'b0000101001010011010 : color = 12'hf01;
15'b0000101001010011011 : color = 12'hf73;
15'b0000101001010011100 : color = 12'he73;
15'b0000101001010011101 : color = 12'hf40;
15'b0000101001010011110 : color = 12'hf00;
15'b0000101001010011111 : color = 12'hf63;
15'b0000101001010100000 : color = 12'he73;
15'b0000101001010100001 : color = 12'he73;
15'b0000101001010100010 : color = 12'he73;
15'b0000101001010100011 : color = 12'he73;
15'b0000101001010100100 : color = 12'he73;
15'b0000101001010100101 : color = 12'he73;
15'b0000101001010100110 : color = 12'he73;
15'b0000101001010100111 : color = 12'he73;
15'b0000101001010101000 : color = 12'he73;
15'b0000101001010101001 : color = 12'he73;
15'b0000101001010101010 : color = 12'he73;
15'b0000101001010101011 : color = 12'he73;
15'b0000101001010101100 : color = 12'he73;
15'b0000101001010101101 : color = 12'he73;
15'b0000101001010101110 : color = 12'he73;
15'b0000101001010101111 : color = 12'he73;
15'b0000101001010110000 : color = 12'he73;
15'b0000101001010110001 : color = 12'he73;
15'b0000101001010110010 : color = 12'he73;
15'b0000101001010110011 : color = 12'he73;
15'b0000101001010110100 : color = 12'he73;
15'b0000101001010110101 : color = 12'he73;
15'b0000101001010110110 : color = 12'he73;
15'b0000101001010110111 : color = 12'he73;
15'b0000101001010111000 : color = 12'he73;
15'b0000101001010111001 : color = 12'he73;
15'b0000101001010111010 : color = 12'he73;
15'b0000101001010111011 : color = 12'he73;
15'b0000101001010111100 : color = 12'he73;
15'b0000101001010111101 : color = 12'he73;
15'b0000101001010111110 : color = 12'he73;
15'b0000101001010111111 : color = 12'he51;
15'b0000101001011000000 : color = 12'hf00;
15'b0000101001011000001 : color = 12'hf63;
15'b0000101001011000010 : color = 12'he73;
15'b0000101001011000011 : color = 12'he73;
15'b0000101001011000100 : color = 12'hf30;
15'b0000101001011000101 : color = 12'hf11;
15'b0000101001011000110 : color = 12'hf73;
15'b0000101001011000111 : color = 12'he73;
15'b0000101001011001000 : color = 12'he73;
15'b0000101001011001001 : color = 12'he73;
15'b0000101001011001010 : color = 12'he61;
15'b0000101001011001011 : color = 12'hf00;
15'b0000101001011001100 : color = 12'hf53;
15'b0000101001011001101 : color = 12'he73;
15'b0000101001011001110 : color = 12'he73;
15'b0000101001011001111 : color = 12'he73;
15'b0000101001011010000 : color = 12'he73;
15'b0000101001011010001 : color = 12'he51;
15'b0000101001011010010 : color = 12'hf00;
15'b0000101001011010011 : color = 12'hf63;
15'b0000101001011010100 : color = 12'he73;
15'b0000101001011010101 : color = 12'he73;
15'b0000101001011010110 : color = 12'he73;
15'b0000101001011010111 : color = 12'he73;
15'b0000101001011011000 : color = 12'he73;
15'b0000101001011011001 : color = 12'he73;
15'b0000101001011011010 : color = 12'he73;
15'b0000101001011011011 : color = 12'he73;
15'b0000101001011011100 : color = 12'he73;
15'b0000101001011011101 : color = 12'he73;
15'b0000101001011011110 : color = 12'he73;
15'b0000101001011011111 : color = 12'he73;
15'b0000101001011100000 : color = 12'he73;
15'b0000101001011100001 : color = 12'he73;
15'b0000101001011100010 : color = 12'he73;
15'b0000101001011100011 : color = 12'he73;
15'b0000101001011100100 : color = 12'he73;
15'b0000101001011100101 : color = 12'he73;
15'b0000101001011100110 : color = 12'he73;
15'b0000101001011100111 : color = 12'he73;
15'b0000101001011101000 : color = 12'he73;
15'b0000101001011101001 : color = 12'he73;
15'b0000101001011101010 : color = 12'he73;
15'b0000101001011101011 : color = 12'he72;
15'b0000101001011101100 : color = 12'hf00;
15'b0000101001011101101 : color = 12'hf11;
15'b0000101001011101110 : color = 12'hf63;
15'b0000101001011101111 : color = 12'he73;
15'b0000101001011110000 : color = 12'he73;
15'b0000101001011110001 : color = 12'he73;
15'b0000101001011110010 : color = 12'he73;
15'b0000101001011110011 : color = 12'he73;
15'b0000101001011110100 : color = 12'he73;
15'b0000101001011110101 : color = 12'he73;
15'b0000101001011110110 : color = 12'he73;
15'b0000101001011110111 : color = 12'he73;
15'b0000101001011111000 : color = 12'he51;
15'b0000101001011111001 : color = 12'hf00;
15'b0000101001011111010 : color = 12'hf53;
15'b0000101001011111011 : color = 12'he73;
15'b0000101001011111100 : color = 12'he73;
15'b0000101001011111101 : color = 12'he73;
15'b0000101001011111110 : color = 12'he73;
15'b0000101001011111111 : color = 12'he73;
15'b0000101001100000000 : color = 12'he73;
15'b0000101001100000001 : color = 12'he73;
15'b0000101001100000010 : color = 12'he73;
15'b0000101001100000011 : color = 12'he73;
15'b0000101001100000100 : color = 12'he73;
15'b0000101001100000101 : color = 12'he73;
15'b0000101001100000110 : color = 12'he73;
15'b0000101001100000111 : color = 12'he73;
15'b0000101001100001000 : color = 12'he73;
15'b0000101001100001001 : color = 12'he73;
15'b0000101001100001010 : color = 12'he73;
15'b0000101001100001011 : color = 12'he73;
15'b0000101001100001100 : color = 12'he73;
15'b0000101001100001101 : color = 12'he73;
15'b0000101001100001110 : color = 12'he73;
15'b0000101001100001111 : color = 12'he73;
15'b0000101001100010000 : color = 12'he73;
15'b0000101001100010001 : color = 12'he73;
15'b0000101001100010010 : color = 12'he73;
15'b0000101001100010011 : color = 12'he73;
15'b0000101001100010100 : color = 12'he73;
15'b0000101001100010101 : color = 12'he73;
15'b0000101001100010110 : color = 12'he73;
15'b0000101001100010111 : color = 12'he73;
15'b0000101001100011000 : color = 12'he73;
15'b0000101001100011001 : color = 12'hf30;
15'b0000101001100011010 : color = 12'hf11;
15'b0000101001100011011 : color = 12'hf73;
15'b0000101001100011100 : color = 12'he73;
15'b0000101001100011101 : color = 12'he73;
15'b0000101001100011110 : color = 12'he73;
15'b0000101001100011111 : color = 12'he73;
15'b0000101001100100000 : color = 12'he73;
15'b0000101001100100001 : color = 12'he73;
15'b0000101001100100010 : color = 12'he73;
15'b0000101001100100011 : color = 12'he73;
15'b0000101001100100100 : color = 12'he72;
15'b0000101001100100101 : color = 12'hf10;
15'b0000101001100100110 : color = 12'hf32;
15'b0000101001100100111 : color = 12'he73;
15'b0000101001100101000 : color = 12'he73;
15'b0000101001100101001 : color = 12'he73;
15'b0000101001100101010 : color = 12'he73;
15'b0000101001100101011 : color = 12'he73;
15'b0000101001100101100 : color = 12'he73;
15'b0000101001100101101 : color = 12'he73;
15'b0000101001100101110 : color = 12'he73;
15'b0000101001100101111 : color = 12'he73;
15'b0000101001100110000 : color = 12'he73;
15'b0000101001100110001 : color = 12'he73;
15'b0000101001100110010 : color = 12'he73;
15'b0000101001100110011 : color = 12'he73;
15'b0000101001100110100 : color = 12'he73;
15'b0000101001100110101 : color = 12'he73;
15'b0000101001100110110 : color = 12'he73;
15'b0000101001100110111 : color = 12'he73;
15'b0000101001100111000 : color = 12'he73;
15'b0000101001100111001 : color = 12'he73;
15'b0000101001100111010 : color = 12'he73;
15'b0000101001100111011 : color = 12'he73;
15'b0000101001100111100 : color = 12'he73;
15'b0000101001100111101 : color = 12'he73;
15'b0000101001100111110 : color = 12'he73;
15'b0000101001100111111 : color = 12'he73;
15'b0000101001101000000 : color = 12'he73;
15'b0000101001101000001 : color = 12'he73;
15'b0000101001101000010 : color = 12'he73;
15'b0000101001101000011 : color = 12'he72;
15'b0000101001101000100 : color = 12'hf10;
15'b0000101001101000101 : color = 12'hf32;
15'b0000101001101000110 : color = 12'he73;
15'b0000101001101000111 : color = 12'he73;
15'b0000101001101001000 : color = 12'he73;
15'b0000101001101001001 : color = 12'he73;
15'b0000101001101001010 : color = 12'he73;
15'b0000101001101001011 : color = 12'he73;
15'b0000101001101001100 : color = 12'he73;
15'b0000101001101001101 : color = 12'he73;
15'b0000101001101001110 : color = 12'he73;
15'b0000101001101001111 : color = 12'he73;
15'b0000101001101010000 : color = 12'hf30;
15'b0000101001101010001 : color = 12'hf32;
15'b0000101001101010010 : color = 12'he73;
15'b0000101001101010011 : color = 12'he73;
15'b0000101001101010100 : color = 12'he73;
15'b0000101001101010101 : color = 12'he73;
15'b0000101001101010110 : color = 12'he73;
15'b0000101001101010111 : color = 12'he73;
15'b0000101001101011000 : color = 12'he73;
15'b0000101001101011001 : color = 12'he73;
15'b0000101001101011010 : color = 12'he73;
15'b0000101001101011011 : color = 12'he73;
15'b0000101001101011100 : color = 12'he73;
15'b0000101001101011101 : color = 12'he73;
15'b0000101001101011110 : color = 12'he73;
15'b0000101001101011111 : color = 12'he73;
15'b0000101001101100000 : color = 12'he73;
15'b0000101001101100001 : color = 12'he73;
15'b0000101001101100010 : color = 12'he73;
15'b0000101001101100011 : color = 12'he73;
15'b0000101001101100100 : color = 12'he73;
15'b0000101001101100101 : color = 12'he73;
15'b0000101001101100110 : color = 12'he73;
15'b0000101001101100111 : color = 12'he73;
15'b0000101001101101000 : color = 12'he73;
15'b0000101001101101001 : color = 12'he73;
15'b0000101001101101010 : color = 12'he73;
15'b0000101001101101011 : color = 12'he73;
15'b0000101001101101100 : color = 12'he73;
15'b0000101001101101101 : color = 12'he73;
15'b0000101001101101110 : color = 12'he73;
15'b0000101001101101111 : color = 12'he73;
15'b0000101001101110000 : color = 12'hf52;
15'b0000101001101110001 : color = 12'hf73;
15'b0000101001101110010 : color = 12'he73;
15'b0000101001101110011 : color = 12'he72;
15'b0000101001101110100 : color = 12'hf63;
15'b0000101001101110101 : color = 12'he73;
15'b0000101001101110110 : color = 12'he73;
15'b0000101001101110111 : color = 12'he73;
15'b0000101001101111000 : color = 12'he51;
15'b0000101001101111001 : color = 12'hf00;
15'b0000101001101111010 : color = 12'hf53;
15'b0000101001101111011 : color = 12'he73;
15'b0000101001101111100 : color = 12'he73;
15'b0000101001101111101 : color = 12'he73;
15'b0000101001101111110 : color = 12'he73;
15'b0000101001101111111 : color = 12'he73;
15'b0000101001110000000 : color = 12'he73;
15'b0000101001110000001 : color = 12'he72;
15'b0000101001110000010 : color = 12'hf11;
15'b0000101001110000011 : color = 12'hf73;
15'b0000101001110000100 : color = 12'he73;
15'b0000101001110000101 : color = 12'he73;
15'b0000101001110000110 : color = 12'he73;
15'b0000101001110000111 : color = 12'he73;
15'b0000101001110001000 : color = 12'he73;
15'b0000101001110001001 : color = 12'he73;
15'b0000101001110001010 : color = 12'he73;
15'b0000101001110001011 : color = 12'he73;
15'b0000101001110001100 : color = 12'he73;
15'b0000101001110001101 : color = 12'he73;
15'b0000101001110001110 : color = 12'he73;
15'b0000101001110001111 : color = 12'he73;
15'b0000101001110010000 : color = 12'he73;
15'b0000101001110010001 : color = 12'he73;
15'b0000101001110010010 : color = 12'he73;
15'b0000101001110010011 : color = 12'he73;
15'b0000101001110010100 : color = 12'he73;
15'b0000101001110010101 : color = 12'he73;
15'b0000101001110010110 : color = 12'he73;
15'b0000101001110010111 : color = 12'he73;
15'b0000101001110011000 : color = 12'he72;
15'b0000101001110011001 : color = 12'hf10;
15'b0000101001110011010 : color = 12'hf32;
15'b0000101001110011011 : color = 12'hf63;
15'b0000101001110011100 : color = 12'he73;
15'b0000101001110011101 : color = 12'he73;
15'b0000101001110011110 : color = 12'he73;
15'b0000101001110011111 : color = 12'he73;
15'b0000101001110100000 : color = 12'he73;
15'b0000101001110100001 : color = 12'he73;
15'b0000101001110100010 : color = 12'he73;
15'b0000101001110100011 : color = 12'he73;
15'b0000101001110100100 : color = 12'he73;
15'b0000101001110100101 : color = 12'he51;
15'b0000101001110100110 : color = 12'hf00;
15'b0000101001110100111 : color = 12'hf53;
15'b0000101001110101000 : color = 12'he73;
15'b0000101001110101001 : color = 12'he73;
15'b0000101001110101010 : color = 12'hf30;
15'b0000101001110101011 : color = 12'hf11;
15'b0000101001110101100 : color = 12'hf73;
15'b0000101001110101101 : color = 12'he73;
15'b0000101001110101110 : color = 12'he73;
15'b0000101001110101111 : color = 12'he73;
15'b0000101001110110000 : color = 12'he73;
15'b0000101001110110001 : color = 12'he73;
15'b0000101001110110010 : color = 12'he73;
15'b0000101001110110011 : color = 12'he73;
15'b0000101001110110100 : color = 12'he73;
15'b0000101001110110101 : color = 12'he73;
15'b0000101001110110110 : color = 12'he73;
15'b0000101001110110111 : color = 12'he73;
15'b0000101001110111000 : color = 12'he73;
15'b0000101001110111001 : color = 12'he73;
15'b0000101001110111010 : color = 12'he73;
15'b0000101001110111011 : color = 12'he73;
15'b0000101001110111100 : color = 12'he73;
15'b0000101001110111101 : color = 12'he73;
15'b0000101001110111110 : color = 12'he73;
15'b0000101001110111111 : color = 12'he73;
15'b0000101001111000000 : color = 12'he73;
15'b0000101001111000001 : color = 12'he73;
15'b0000101001000000000 : color = 12'he73;
15'b0000101001000000001 : color = 12'he73;
15'b0000101001000000010 : color = 12'he73;
15'b0000101001000000011 : color = 12'he73;
15'b0000101001000000100 : color = 12'he73;
15'b0000101001000000101 : color = 12'he73;
15'b0000101001000000110 : color = 12'he73;
15'b0000101001000000111 : color = 12'he73;
15'b0000101001000001000 : color = 12'he73;
15'b0000101001000001001 : color = 12'he73;
15'b0000101001000001010 : color = 12'he73;
15'b0000101001000001011 : color = 12'he72;
15'b0000101001000001100 : color = 12'hf00;
15'b0000101001000001101 : color = 12'hf63;
15'b0000101001000001110 : color = 12'he73;
15'b0000101001000001111 : color = 12'he73;
15'b0000101001000010000 : color = 12'he51;
15'b0000101001000010001 : color = 12'hf00;
15'b0000101001000010010 : color = 12'hf01;
15'b0000101001000010011 : color = 12'hf73;
15'b0000101001000010100 : color = 12'he73;
15'b0000101001000010101 : color = 12'he73;
15'b0000101001000010110 : color = 12'he72;
15'b0000101001000010111 : color = 12'hf10;
15'b0000101001000011000 : color = 12'hf32;
15'b0000101001000011001 : color = 12'he73;
15'b0000101001000011010 : color = 12'he73;
15'b0000101001000011011 : color = 12'he61;
15'b0000101001000011100 : color = 12'hf01;
15'b0000101001000011101 : color = 12'hf73;
15'b0000101001000011110 : color = 12'he73;
15'b0000101001000011111 : color = 12'he73;
15'b0000101001000100000 : color = 12'he73;
15'b0000101001000100001 : color = 12'he73;
15'b0000101001000100010 : color = 12'he73;
15'b0000101001000100011 : color = 12'he73;
15'b0000101001000100100 : color = 12'he73;
15'b0000101001000100101 : color = 12'he73;
15'b0000101001000100110 : color = 12'he73;
15'b0000101001000100111 : color = 12'he73;
15'b0000101001000101000 : color = 12'he73;
15'b0000101001000101001 : color = 12'he73;
15'b0000101001000101010 : color = 12'he73;
15'b0000101001000101011 : color = 12'he73;
15'b0000101001000101100 : color = 12'he73;
15'b0000101001000101101 : color = 12'he73;
15'b0000101001000101110 : color = 12'he73;
15'b0000101001000101111 : color = 12'he73;
15'b0000101001000110000 : color = 12'he73;
15'b0000101001000110001 : color = 12'he73;
15'b0000101001000110010 : color = 12'he73;
15'b0000101001000110011 : color = 12'he73;
15'b0000101001000110100 : color = 12'he73;
15'b0000101001000110101 : color = 12'he73;
15'b0000101001000110110 : color = 12'he73;
15'b0000101001000110111 : color = 12'he73;
15'b0000101001000111000 : color = 12'he51;
15'b0000101001000111001 : color = 12'hf00;
15'b0000101001000111010 : color = 12'hf63;
15'b0000101001000111011 : color = 12'he73;
15'b0000101001000111100 : color = 12'he73;
15'b0000101001000111101 : color = 12'he72;
15'b0000101001000111110 : color = 12'hf10;
15'b0000101001000111111 : color = 12'hf42;
15'b0000101001001000000 : color = 12'he73;
15'b0000101001001000001 : color = 12'he73;
15'b0000101001001000010 : color = 12'he73;
15'b0000101001001000011 : color = 12'he73;
15'b0000101001001000100 : color = 12'he72;
15'b0000101001001000101 : color = 12'hf10;
15'b0000101001001000110 : color = 12'hf32;
15'b0000101001001000111 : color = 12'he73;
15'b0000101001001001000 : color = 12'he73;
15'b0000101001001001001 : color = 12'he62;
15'b0000101001001001010 : color = 12'hf00;
15'b0000101001001001011 : color = 12'hf00;
15'b0000101001001001100 : color = 12'hf63;
15'b0000101001001001101 : color = 12'he73;
15'b0000101001001001110 : color = 12'he73;
15'b0000101001001001111 : color = 12'he73;
15'b0000101001001010000 : color = 12'he73;
15'b0000101001001010001 : color = 12'he73;
15'b0000101001001010010 : color = 12'he73;
15'b0000101001001010011 : color = 12'he73;
15'b0000101001001010100 : color = 12'he73;
15'b0000101001001010101 : color = 12'he73;
15'b0000101001001010110 : color = 12'he73;
15'b0000101001001010111 : color = 12'he73;
15'b0000101001001011000 : color = 12'he73;
15'b0000101001001011001 : color = 12'he73;
15'b0000101001001011010 : color = 12'he73;
15'b0000101001001011011 : color = 12'he73;
15'b0000101001001011100 : color = 12'he73;
15'b0000101001001011101 : color = 12'he73;
15'b0000101001001011110 : color = 12'he73;
15'b0000101001001011111 : color = 12'he73;
15'b0000101001001100000 : color = 12'he73;
15'b0000101001001100001 : color = 12'he73;
15'b0000101001001100010 : color = 12'he73;
15'b0000101001001100011 : color = 12'he73;
15'b0000101001001100100 : color = 12'he73;
15'b0000101001001100101 : color = 12'he73;
15'b0000101001001100110 : color = 12'he73;
15'b0000101001001100111 : color = 12'he73;
15'b0000101001001101000 : color = 12'hf40;
15'b0000101001001101001 : color = 12'hf00;
15'b0000101001001101010 : color = 12'hf53;
15'b0000101001001101011 : color = 12'he73;
15'b0000101001001101100 : color = 12'he51;
15'b0000101001001101101 : color = 12'hf00;
15'b0000101001001101110 : color = 12'hf53;
15'b0000101001001101111 : color = 12'he73;
15'b0000101001001110000 : color = 12'he72;
15'b0000101001001110001 : color = 12'hf10;
15'b0000101001001110010 : color = 12'hf32;
15'b0000101001001110011 : color = 12'hf73;
15'b0000101001001110100 : color = 12'he73;
15'b0000101001001110101 : color = 12'he73;
15'b0000101001001110110 : color = 12'he73;
15'b0000101001001110111 : color = 12'he73;
15'b0000101001001111000 : color = 12'he73;
15'b0000101001001111001 : color = 12'he73;
15'b0000101001001111010 : color = 12'he73;
15'b0000101001001111011 : color = 12'he73;
15'b0000101001001111100 : color = 12'he73;
15'b0000101001001111101 : color = 12'he73;
15'b0000101001001111110 : color = 12'he73;
15'b0000101001001111111 : color = 12'he73;
15'b0000101001010000000 : color = 12'he73;
15'b0000101001010000001 : color = 12'he73;
15'b0000101001010000010 : color = 12'he73;
15'b0000101001010000011 : color = 12'he73;
15'b0000101001010000100 : color = 12'he73;
15'b0000101001010000101 : color = 12'he73;
15'b0000101001010000110 : color = 12'he73;
15'b0000101001010000111 : color = 12'he73;
15'b0000101001010001000 : color = 12'he73;
15'b0000101001010001001 : color = 12'he73;
15'b0000101001010001010 : color = 12'he73;
15'b0000101001010001011 : color = 12'he73;
15'b0000101001010001100 : color = 12'he73;
15'b0000101001010001101 : color = 12'he73;
15'b0000101001010001110 : color = 12'he73;
15'b0000101001010001111 : color = 12'he73;
15'b0000101001010010000 : color = 12'he73;
15'b0000101001010010001 : color = 12'he73;
15'b0000101001010010010 : color = 12'he73;
15'b0000101001010010011 : color = 12'he72;
15'b0000101001010010100 : color = 12'hf00;
15'b0000101001010010101 : color = 12'hf42;
15'b0000101001010010110 : color = 12'he73;
15'b0000101001010010111 : color = 12'he73;
15'b0000101001010011000 : color = 12'he73;
15'b0000101001010011001 : color = 12'he73;
15'b0000101001010011010 : color = 12'he73;
15'b0000101001010011011 : color = 12'he73;
15'b0000101001010011100 : color = 12'he73;
15'b0000101001010011101 : color = 12'he72;
15'b0000101001010011110 : color = 12'hf10;
15'b0000101001010011111 : color = 12'hf32;
15'b0000101001010100000 : color = 12'he73;
15'b0000101001010100001 : color = 12'he73;
15'b0000101001010100010 : color = 12'he73;
15'b0000101001010100011 : color = 12'hf40;
15'b0000101001010100100 : color = 12'hf01;
15'b0000101001010100101 : color = 12'hf73;
15'b0000101001010100110 : color = 12'he73;
15'b0000101001010100111 : color = 12'he73;
15'b0000101001010101000 : color = 12'he73;
15'b0000101001010101001 : color = 12'he73;
15'b0000101001010101010 : color = 12'he73;
15'b0000101001010101011 : color = 12'he73;
15'b0000101001010101100 : color = 12'he73;
15'b0000101001010101101 : color = 12'he73;
15'b0000101001010101110 : color = 12'he73;
15'b0000101001010101111 : color = 12'he73;
15'b0000101001010110000 : color = 12'he73;
15'b0000101001010110001 : color = 12'he73;
15'b0000101001010110010 : color = 12'he73;
15'b0000101001010110011 : color = 12'he73;
15'b0000101001010110100 : color = 12'he73;
15'b0000101001010110101 : color = 12'he73;
15'b0000101001010110110 : color = 12'he73;
15'b0000101001010110111 : color = 12'he73;
15'b0000101001010111000 : color = 12'he73;
15'b0000101001010111001 : color = 12'he73;
15'b0000101001010111010 : color = 12'he73;
15'b0000101001010111011 : color = 12'he73;
15'b0000101001010111100 : color = 12'he73;
15'b0000101001010111101 : color = 12'he73;
15'b0000101001010111110 : color = 12'he73;
15'b0000101001010111111 : color = 12'he73;
15'b0000101001011000000 : color = 12'he73;
15'b0000101001011000001 : color = 12'he73;
15'b0000101001011000010 : color = 12'he72;
15'b0000101001011000011 : color = 12'hf10;
15'b0000101001011000100 : color = 12'hf32;
15'b0000101001011000101 : color = 12'hf61;
15'b0000101001011000110 : color = 12'hf00;
15'b0000101001011000111 : color = 12'hf42;
15'b0000101001011001000 : color = 12'he73;
15'b0000101001011001001 : color = 12'he73;
15'b0000101001011001010 : color = 12'he73;
15'b0000101001011001011 : color = 12'he73;
15'b0000101001011001100 : color = 12'he73;
15'b0000101001011001101 : color = 12'he73;
15'b0000101001011001110 : color = 12'he73;
15'b0000101001011001111 : color = 12'he73;
15'b0000101001011010000 : color = 12'he73;
15'b0000101001011010001 : color = 12'he73;
15'b0000101001011010010 : color = 12'he73;
15'b0000101001011010011 : color = 12'he73;
15'b0000101001011010100 : color = 12'he73;
15'b0000101001011010101 : color = 12'he73;
15'b0000101001011010110 : color = 12'he73;
15'b0000101001011010111 : color = 12'he73;
15'b0000101001011011000 : color = 12'he73;
15'b0000101001011011001 : color = 12'he73;
15'b0000101001011011010 : color = 12'he73;
15'b0000101001011011011 : color = 12'he73;
15'b0000101001011011100 : color = 12'he73;
15'b0000101001011011101 : color = 12'he73;
15'b0000101001011011110 : color = 12'he73;
15'b0000101001011011111 : color = 12'he73;
15'b0000101001011100000 : color = 12'he73;
15'b0000101001011100001 : color = 12'he73;
15'b0000101001011100010 : color = 12'he73;
15'b0000101001011100011 : color = 12'he73;
15'b0000101001011100100 : color = 12'he73;
15'b0000101001011100101 : color = 12'he73;
15'b0000101001011100110 : color = 12'he73;
15'b0000101001011100111 : color = 12'he73;
15'b0000101001011101000 : color = 12'he51;
15'b0000101001011101001 : color = 12'hf00;
15'b0000101001011101010 : color = 12'hf63;
15'b0000101001011101011 : color = 12'he73;
15'b0000101001011101100 : color = 12'he73;
15'b0000101001011101101 : color = 12'hf30;
15'b0000101001011101110 : color = 12'hf11;
15'b0000101001011101111 : color = 12'hf73;
15'b0000101001011110000 : color = 12'he73;
15'b0000101001011110001 : color = 12'he73;
15'b0000101001011110010 : color = 12'he73;
15'b0000101001011110011 : color = 12'he61;
15'b0000101001011110100 : color = 12'hf00;
15'b0000101001011110101 : color = 12'hf53;
15'b0000101001011110110 : color = 12'he73;
15'b0000101001011110111 : color = 12'he73;
15'b0000101001011111000 : color = 12'he73;
15'b0000101001011111001 : color = 12'he73;
15'b0000101001011111010 : color = 12'he51;
15'b0000101001011111011 : color = 12'hf00;
15'b0000101001011111100 : color = 12'hf63;
15'b0000101001011111101 : color = 12'he73;
15'b0000101001011111110 : color = 12'he73;
15'b0000101001011111111 : color = 12'he73;
15'b0000101001100000000 : color = 12'he73;
15'b0000101001100000001 : color = 12'he73;
15'b0000101001100000010 : color = 12'he73;
15'b0000101001100000011 : color = 12'he73;
15'b0000101001100000100 : color = 12'he73;
15'b0000101001100000101 : color = 12'he73;
15'b0000101001100000110 : color = 12'he73;
15'b0000101001100000111 : color = 12'he73;
15'b0000101001100001000 : color = 12'he73;
15'b0000101001100001001 : color = 12'he73;
15'b0000101001100001010 : color = 12'he73;
15'b0000101001100001011 : color = 12'he73;
15'b0000101001100001100 : color = 12'he73;
15'b0000101001100001101 : color = 12'he73;
15'b0000101001100001110 : color = 12'he73;
15'b0000101001100001111 : color = 12'he73;
15'b0000101001100010000 : color = 12'he73;
15'b0000101001100010001 : color = 12'he73;
15'b0000101001100010010 : color = 12'he73;
15'b0000101001100010011 : color = 12'he73;
15'b0000101001100010100 : color = 12'he61;
15'b0000101001100010101 : color = 12'hf00;
15'b0000101001100010110 : color = 12'hf52;
15'b0000101001100010111 : color = 12'hf30;
15'b0000101001100011000 : color = 12'hf32;
15'b0000101001100011001 : color = 12'hf73;
15'b0000101001100011010 : color = 12'he73;
15'b0000101001100011011 : color = 12'he73;
15'b0000101001100011100 : color = 12'he73;
15'b0000101001100011101 : color = 12'he73;
15'b0000101001100011110 : color = 12'he73;
15'b0000101001100011111 : color = 12'he73;
15'b0000101001100100000 : color = 12'he73;
15'b0000101001100100001 : color = 12'he51;
15'b0000101001100100010 : color = 12'hf00;
15'b0000101001100100011 : color = 12'hf53;
15'b0000101001100100100 : color = 12'he73;
15'b0000101001100100101 : color = 12'he73;
15'b0000101001100100110 : color = 12'he73;
15'b0000101001100100111 : color = 12'he73;
15'b0000101001100101000 : color = 12'he73;
15'b0000101001100101001 : color = 12'he73;
15'b0000101001100101010 : color = 12'he73;
15'b0000101001100101011 : color = 12'he73;
15'b0000101001100101100 : color = 12'he73;
15'b0000101001100101101 : color = 12'he73;
15'b0000101001100101110 : color = 12'he73;
15'b0000101001100101111 : color = 12'he73;
15'b0000101001100110000 : color = 12'he73;
15'b0000101001100110001 : color = 12'he73;
15'b0000101001100110010 : color = 12'he73;
15'b0000101001100110011 : color = 12'he73;
15'b0000101001100110100 : color = 12'he73;
15'b0000101001100110101 : color = 12'he73;
15'b0000101001100110110 : color = 12'he73;
15'b0000101001100110111 : color = 12'he73;
15'b0000101001100111000 : color = 12'he73;
15'b0000101001100111001 : color = 12'he73;
15'b0000101001100111010 : color = 12'he73;
15'b0000101001100111011 : color = 12'he73;
15'b0000101001100111100 : color = 12'he73;
15'b0000101001100111101 : color = 12'he73;
15'b0000101001100111110 : color = 12'he73;
15'b0000101001100111111 : color = 12'he73;
15'b0000101001101000000 : color = 12'he73;
15'b0000101001101000001 : color = 12'he73;
15'b0000101001101000010 : color = 12'hf30;
15'b0000101001101000011 : color = 12'hf11;
15'b0000101001101000100 : color = 12'hf73;
15'b0000101001101000101 : color = 12'he73;
15'b0000101001101000110 : color = 12'he73;
15'b0000101001101000111 : color = 12'he73;
15'b0000101001101001000 : color = 12'he73;
15'b0000101001101001001 : color = 12'he73;
15'b0000101001101001010 : color = 12'he73;
15'b0000101001101001011 : color = 12'he73;
15'b0000101001101001100 : color = 12'he73;
15'b0000101001101001101 : color = 12'he73;
15'b0000101001101001110 : color = 12'he73;
15'b0000101001101001111 : color = 12'he73;
15'b0000101001101010000 : color = 12'he73;
15'b0000101001101010001 : color = 12'he73;
15'b0000101001101010010 : color = 12'he73;
15'b0000101001101010011 : color = 12'he73;
15'b0000101001101010100 : color = 12'he73;
15'b0000101001101010101 : color = 12'he73;
15'b0000101001101010110 : color = 12'he73;
15'b0000101001101010111 : color = 12'he73;
15'b0000101001101011000 : color = 12'he73;
15'b0000101001101011001 : color = 12'he73;
15'b0000101001101011010 : color = 12'he73;
15'b0000101001101011011 : color = 12'he73;
15'b0000101001101011100 : color = 12'he73;
15'b0000101001101011101 : color = 12'he73;
15'b0000101001101011110 : color = 12'he73;
15'b0000101001101011111 : color = 12'he73;
15'b0000101001101100000 : color = 12'he73;
15'b0000101001101100001 : color = 12'he73;
15'b0000101001101100010 : color = 12'he73;
15'b0000101001101100011 : color = 12'he73;
15'b0000101001101100100 : color = 12'he73;
15'b0000101001101100101 : color = 12'he73;
15'b0000101001101100110 : color = 12'he73;
15'b0000101001101100111 : color = 12'he73;
15'b0000101001101101000 : color = 12'he73;
15'b0000101001101101001 : color = 12'he73;
15'b0000101001101101010 : color = 12'he73;
15'b0000101001101101011 : color = 12'he73;
15'b0000101001101101100 : color = 12'he72;
15'b0000101001101101101 : color = 12'hf10;
15'b0000101001101101110 : color = 12'hf32;
15'b0000101001101101111 : color = 12'he73;
15'b0000101001101110000 : color = 12'he73;
15'b0000101001101110001 : color = 12'he73;
15'b0000101001101110010 : color = 12'he62;
15'b0000101001101110011 : color = 12'hf63;
15'b0000101001101110100 : color = 12'he73;
15'b0000101001101110101 : color = 12'he73;
15'b0000101001101110110 : color = 12'he73;
15'b0000101001101110111 : color = 12'he73;
15'b0000101001101111000 : color = 12'he73;
15'b0000101001101111001 : color = 12'hf30;
15'b0000101001101111010 : color = 12'hf32;
15'b0000101001101111011 : color = 12'he73;
15'b0000101001101111100 : color = 12'he73;
15'b0000101001101111101 : color = 12'he73;
15'b0000101001101111110 : color = 12'he61;
15'b0000101001101111111 : color = 12'hf11;
15'b0000101001110000000 : color = 12'hf73;
15'b0000101001110000001 : color = 12'he73;
15'b0000101001110000010 : color = 12'he73;
15'b0000101001110000011 : color = 12'he73;
15'b0000101001110000100 : color = 12'he73;
15'b0000101001110000101 : color = 12'he73;
15'b0000101001110000110 : color = 12'he73;
15'b0000101001110000111 : color = 12'he73;
15'b0000101001110001000 : color = 12'he73;
15'b0000101001110001001 : color = 12'he73;
15'b0000101001110001010 : color = 12'he73;
15'b0000101001110001011 : color = 12'he73;
15'b0000101001110001100 : color = 12'he73;
15'b0000101001110001101 : color = 12'he73;
15'b0000101001110001110 : color = 12'he73;
15'b0000101001110001111 : color = 12'he73;
15'b0000101001110010000 : color = 12'he73;
15'b0000101001110010001 : color = 12'he73;
15'b0000101001110010010 : color = 12'he73;
15'b0000101001110010011 : color = 12'he73;
15'b0000101001110010100 : color = 12'he73;
15'b0000101001110010101 : color = 12'he73;
15'b0000101001110010110 : color = 12'he73;
15'b0000101001110010111 : color = 12'he73;
15'b0000101001110011000 : color = 12'he73;
15'b0000101001110011001 : color = 12'he73;
15'b0000101001110011010 : color = 12'he73;
15'b0000101001110011011 : color = 12'he73;
15'b0000101001110011100 : color = 12'hf40;
15'b0000101001110011101 : color = 12'hf00;
15'b0000101001110011110 : color = 12'hf63;
15'b0000101001110011111 : color = 12'he73;
15'b0000101001110100000 : color = 12'he73;
15'b0000101001110100001 : color = 12'he51;
15'b0000101001110100010 : color = 12'hf00;
15'b0000101001110100011 : color = 12'hf53;
15'b0000101001110100100 : color = 12'he72;
15'b0000101001110100101 : color = 12'hf31;
15'b0000101001110100110 : color = 12'hf52;
15'b0000101001110100111 : color = 12'hf73;
15'b0000101001110101000 : color = 12'he73;
15'b0000101001110101001 : color = 12'he73;
15'b0000101001110101010 : color = 12'he73;
15'b0000101001110101011 : color = 12'he73;
15'b0000101001110101100 : color = 12'he73;
15'b0000101001110101101 : color = 12'he73;
15'b0000101001110101110 : color = 12'he73;
15'b0000101001110101111 : color = 12'he73;
15'b0000101001110110000 : color = 12'he73;
15'b0000101001110110001 : color = 12'he73;
15'b0000101001110110010 : color = 12'he73;
15'b0000101001110110011 : color = 12'he73;
15'b0000101001110110100 : color = 12'he73;
15'b0000101001110110101 : color = 12'he73;
15'b0000101001110110110 : color = 12'he73;
15'b0000101001110110111 : color = 12'he73;
15'b0000101001110111000 : color = 12'he73;
15'b0000101001110111001 : color = 12'he73;
15'b0000101001110111010 : color = 12'he73;
15'b0000101001110111011 : color = 12'he73;
15'b0000101001110111100 : color = 12'he73;
15'b0000101001110111101 : color = 12'he73;
15'b0000101001110111110 : color = 12'he73;
15'b0000101001110111111 : color = 12'he73;
15'b0000101001111000000 : color = 12'he73;
15'b0000101001111000001 : color = 12'he73;
15'b0000101001111000010 : color = 12'he73;
15'b0000101001111000011 : color = 12'he73;
15'b0000101001111000100 : color = 12'he73;
15'b0000101001111000101 : color = 12'he73;
15'b0000101001111000110 : color = 12'he73;
15'b0000101001111000111 : color = 12'he73;
15'b0000101001111001000 : color = 12'he73;
15'b0000101001111001001 : color = 12'he73;
15'b0000101001111001010 : color = 12'he73;
15'b0000101001111001011 : color = 12'he73;
15'b0000101001111001100 : color = 12'he73;
15'b0000101001111001101 : color = 12'he73;
15'b0000101001111001110 : color = 12'he51;
15'b0000101001111001111 : color = 12'hf00;
15'b0000101001111010000 : color = 12'hf63;
15'b0000101001111010001 : color = 12'he73;
15'b0000101001111010010 : color = 12'he73;
15'b0000101001111010011 : color = 12'hf30;
15'b0000101001111010100 : color = 12'hf11;
15'b0000101001111010101 : color = 12'hf73;
15'b0000101001111010110 : color = 12'he73;
15'b0000101001111010111 : color = 12'he73;
15'b0000101001111011000 : color = 12'he73;
15'b0000101001111011001 : color = 12'he73;
15'b0000101001111011010 : color = 12'he73;
15'b0000101001111011011 : color = 12'he73;
15'b0000101001111011100 : color = 12'he73;
15'b0000101001111011101 : color = 12'he73;
15'b0000101001111011110 : color = 12'he73;
15'b0000101001111011111 : color = 12'he73;
15'b0000101001111100000 : color = 12'he73;
15'b0000101001111100001 : color = 12'he73;
15'b0000101001111100010 : color = 12'he73;
15'b0000101001111100011 : color = 12'he73;
15'b0000101001111100100 : color = 12'he73;
15'b0000101001111100101 : color = 12'he73;
15'b0000101001111100110 : color = 12'he73;
15'b0000101001111100111 : color = 12'he73;
15'b0000101001111101000 : color = 12'he73;
15'b0000101001111101001 : color = 12'he73;
15'b0000101001111101010 : color = 12'he73;
15'b0000101001000101001 : color = 12'he73;
15'b0000101001000101010 : color = 12'he73;
15'b0000101001000101011 : color = 12'he73;
15'b0000101001000101100 : color = 12'he73;
15'b0000101001000101101 : color = 12'he73;
15'b0000101001000101110 : color = 12'he73;
15'b0000101001000101111 : color = 12'he73;
15'b0000101001000110000 : color = 12'he73;
15'b0000101001000110001 : color = 12'he73;
15'b0000101001000110010 : color = 12'he73;
15'b0000101001000110011 : color = 12'he73;
15'b0000101001000110100 : color = 12'hf30;
15'b0000101001000110101 : color = 12'hf42;
15'b0000101001000110110 : color = 12'he73;
15'b0000101001000110111 : color = 12'he73;
15'b0000101001000111000 : color = 12'he73;
15'b0000101001000111001 : color = 12'he72;
15'b0000101001000111010 : color = 12'hf10;
15'b0000101001000111011 : color = 12'hf00;
15'b0000101001000111100 : color = 12'hf53;
15'b0000101001000111101 : color = 12'he73;
15'b0000101001000111110 : color = 12'he73;
15'b0000101001000111111 : color = 12'hf40;
15'b0000101001001000000 : color = 12'hf00;
15'b0000101001001000001 : color = 12'hf63;
15'b0000101001001000010 : color = 12'he73;
15'b0000101001001000011 : color = 12'he73;
15'b0000101001001000100 : color = 12'he72;
15'b0000101001001000101 : color = 12'hf10;
15'b0000101001001000110 : color = 12'hf42;
15'b0000101001001000111 : color = 12'he73;
15'b0000101001001001000 : color = 12'he73;
15'b0000101001001001001 : color = 12'he73;
15'b0000101001001001010 : color = 12'he73;
15'b0000101001001001011 : color = 12'he73;
15'b0000101001001001100 : color = 12'he73;
15'b0000101001001001101 : color = 12'he73;
15'b0000101001001001110 : color = 12'he73;
15'b0000101001001001111 : color = 12'he73;
15'b0000101001001010000 : color = 12'he73;
15'b0000101001001010001 : color = 12'he73;
15'b0000101001001010010 : color = 12'he73;
15'b0000101001001010011 : color = 12'he73;
15'b0000101001001010100 : color = 12'he73;
15'b0000101001001010101 : color = 12'he73;
15'b0000101001001010110 : color = 12'he73;
15'b0000101001001010111 : color = 12'he73;
15'b0000101001001011000 : color = 12'he73;
15'b0000101001001011001 : color = 12'he73;
15'b0000101001001011010 : color = 12'he73;
15'b0000101001001011011 : color = 12'he73;
15'b0000101001001011100 : color = 12'he73;
15'b0000101001001011101 : color = 12'he73;
15'b0000101001001011110 : color = 12'he73;
15'b0000101001001011111 : color = 12'he73;
15'b0000101001001100000 : color = 12'he73;
15'b0000101001001100001 : color = 12'he51;
15'b0000101001001100010 : color = 12'hf00;
15'b0000101001001100011 : color = 12'hf63;
15'b0000101001001100100 : color = 12'he73;
15'b0000101001001100101 : color = 12'he73;
15'b0000101001001100110 : color = 12'he73;
15'b0000101001001100111 : color = 12'he73;
15'b0000101001001101000 : color = 12'he73;
15'b0000101001001101001 : color = 12'he73;
15'b0000101001001101010 : color = 12'he73;
15'b0000101001001101011 : color = 12'he73;
15'b0000101001001101100 : color = 12'he73;
15'b0000101001001101101 : color = 12'he72;
15'b0000101001001101110 : color = 12'hf10;
15'b0000101001001101111 : color = 12'hf32;
15'b0000101001001110000 : color = 12'he73;
15'b0000101001001110001 : color = 12'he73;
15'b0000101001001110010 : color = 12'he73;
15'b0000101001001110011 : color = 12'hf51;
15'b0000101001001110100 : color = 12'hf63;
15'b0000101001001110101 : color = 12'he73;
15'b0000101001001110110 : color = 12'he73;
15'b0000101001001110111 : color = 12'he73;
15'b0000101001001111000 : color = 12'he73;
15'b0000101001001111001 : color = 12'he73;
15'b0000101001001111010 : color = 12'he73;
15'b0000101001001111011 : color = 12'he73;
15'b0000101001001111100 : color = 12'he73;
15'b0000101001001111101 : color = 12'he73;
15'b0000101001001111110 : color = 12'he73;
15'b0000101001001111111 : color = 12'he73;
15'b0000101001010000000 : color = 12'he73;
15'b0000101001010000001 : color = 12'he73;
15'b0000101001010000010 : color = 12'he73;
15'b0000101001010000011 : color = 12'he73;
15'b0000101001010000100 : color = 12'he73;
15'b0000101001010000101 : color = 12'he73;
15'b0000101001010000110 : color = 12'he73;
15'b0000101001010000111 : color = 12'he73;
15'b0000101001010001000 : color = 12'he73;
15'b0000101001010001001 : color = 12'he73;
15'b0000101001010001010 : color = 12'he73;
15'b0000101001010001011 : color = 12'he73;
15'b0000101001010001100 : color = 12'he73;
15'b0000101001010001101 : color = 12'he73;
15'b0000101001010001110 : color = 12'he73;
15'b0000101001010001111 : color = 12'he73;
15'b0000101001010010000 : color = 12'he51;
15'b0000101001010010001 : color = 12'hf00;
15'b0000101001010010010 : color = 12'hf42;
15'b0000101001010010011 : color = 12'he73;
15'b0000101001010010100 : color = 12'he73;
15'b0000101001010010101 : color = 12'hf40;
15'b0000101001010010110 : color = 12'hf00;
15'b0000101001010010111 : color = 12'hf53;
15'b0000101001010011000 : color = 12'he73;
15'b0000101001010011001 : color = 12'he73;
15'b0000101001010011010 : color = 12'he72;
15'b0000101001010011011 : color = 12'hf00;
15'b0000101001010011100 : color = 12'hf11;
15'b0000101001010011101 : color = 12'hf73;
15'b0000101001010011110 : color = 12'he73;
15'b0000101001010011111 : color = 12'he73;
15'b0000101001010100000 : color = 12'he73;
15'b0000101001010100001 : color = 12'he73;
15'b0000101001010100010 : color = 12'he73;
15'b0000101001010100011 : color = 12'he73;
15'b0000101001010100100 : color = 12'he73;
15'b0000101001010100101 : color = 12'he73;
15'b0000101001010100110 : color = 12'he73;
15'b0000101001010100111 : color = 12'he73;
15'b0000101001010101000 : color = 12'he73;
15'b0000101001010101001 : color = 12'he73;
15'b0000101001010101010 : color = 12'he73;
15'b0000101001010101011 : color = 12'he73;
15'b0000101001010101100 : color = 12'he73;
15'b0000101001010101101 : color = 12'he73;
15'b0000101001010101110 : color = 12'he73;
15'b0000101001010101111 : color = 12'he73;
15'b0000101001010110000 : color = 12'he73;
15'b0000101001010110001 : color = 12'he73;
15'b0000101001010110010 : color = 12'he73;
15'b0000101001010110011 : color = 12'he73;
15'b0000101001010110100 : color = 12'he73;
15'b0000101001010110101 : color = 12'he73;
15'b0000101001010110110 : color = 12'he73;
15'b0000101001010110111 : color = 12'he73;
15'b0000101001010111000 : color = 12'he73;
15'b0000101001010111001 : color = 12'he73;
15'b0000101001010111010 : color = 12'he73;
15'b0000101001010111011 : color = 12'he73;
15'b0000101001010111100 : color = 12'he72;
15'b0000101001010111101 : color = 12'hf00;
15'b0000101001010111110 : color = 12'hf42;
15'b0000101001010111111 : color = 12'he73;
15'b0000101001011000000 : color = 12'he73;
15'b0000101001011000001 : color = 12'he73;
15'b0000101001011000010 : color = 12'he73;
15'b0000101001011000011 : color = 12'he73;
15'b0000101001011000100 : color = 12'he73;
15'b0000101001011000101 : color = 12'he73;
15'b0000101001011000110 : color = 12'he72;
15'b0000101001011000111 : color = 12'hf00;
15'b0000101001011001000 : color = 12'hf32;
15'b0000101001011001001 : color = 12'he73;
15'b0000101001011001010 : color = 12'he73;
15'b0000101001011001011 : color = 12'he73;
15'b0000101001011001100 : color = 12'hf40;
15'b0000101001011001101 : color = 12'hf01;
15'b0000101001011001110 : color = 12'hf73;
15'b0000101001011001111 : color = 12'he73;
15'b0000101001011010000 : color = 12'he73;
15'b0000101001011010001 : color = 12'he73;
15'b0000101001011010010 : color = 12'he73;
15'b0000101001011010011 : color = 12'he73;
15'b0000101001011010100 : color = 12'he73;
15'b0000101001011010101 : color = 12'he73;
15'b0000101001011010110 : color = 12'he73;
15'b0000101001011010111 : color = 12'he73;
15'b0000101001011011000 : color = 12'he73;
15'b0000101001011011001 : color = 12'he73;
15'b0000101001011011010 : color = 12'he73;
15'b0000101001011011011 : color = 12'he73;
15'b0000101001011011100 : color = 12'he73;
15'b0000101001011011101 : color = 12'he73;
15'b0000101001011011110 : color = 12'he73;
15'b0000101001011011111 : color = 12'he73;
15'b0000101001011100000 : color = 12'he73;
15'b0000101001011100001 : color = 12'he73;
15'b0000101001011100010 : color = 12'he73;
15'b0000101001011100011 : color = 12'he73;
15'b0000101001011100100 : color = 12'he73;
15'b0000101001011100101 : color = 12'he73;
15'b0000101001011100110 : color = 12'he73;
15'b0000101001011100111 : color = 12'he73;
15'b0000101001011101000 : color = 12'he73;
15'b0000101001011101001 : color = 12'he73;
15'b0000101001011101010 : color = 12'he73;
15'b0000101001011101011 : color = 12'he73;
15'b0000101001011101100 : color = 12'he61;
15'b0000101001011101101 : color = 12'hf00;
15'b0000101001011101110 : color = 12'hf00;
15'b0000101001011101111 : color = 12'hf11;
15'b0000101001011110000 : color = 12'hf73;
15'b0000101001011110001 : color = 12'he73;
15'b0000101001011110010 : color = 12'he73;
15'b0000101001011110011 : color = 12'he73;
15'b0000101001011110100 : color = 12'he73;
15'b0000101001011110101 : color = 12'he73;
15'b0000101001011110110 : color = 12'he73;
15'b0000101001011110111 : color = 12'he73;
15'b0000101001011111000 : color = 12'he73;
15'b0000101001011111001 : color = 12'he73;
15'b0000101001011111010 : color = 12'he73;
15'b0000101001011111011 : color = 12'he73;
15'b0000101001011111100 : color = 12'he73;
15'b0000101001011111101 : color = 12'he73;
15'b0000101001011111110 : color = 12'he73;
15'b0000101001011111111 : color = 12'he73;
15'b0000101001100000000 : color = 12'he73;
15'b0000101001100000001 : color = 12'he73;
15'b0000101001100000010 : color = 12'he73;
15'b0000101001100000011 : color = 12'he73;
15'b0000101001100000100 : color = 12'he73;
15'b0000101001100000101 : color = 12'he73;
15'b0000101001100000110 : color = 12'he73;
15'b0000101001100000111 : color = 12'he73;
15'b0000101001100001000 : color = 12'he73;
15'b0000101001100001001 : color = 12'he73;
15'b0000101001100001010 : color = 12'he73;
15'b0000101001100001011 : color = 12'he73;
15'b0000101001100001100 : color = 12'he73;
15'b0000101001100001101 : color = 12'he73;
15'b0000101001100001110 : color = 12'he73;
15'b0000101001100001111 : color = 12'he73;
15'b0000101001100010000 : color = 12'he73;
15'b0000101001100010001 : color = 12'he51;
15'b0000101001100010010 : color = 12'hf00;
15'b0000101001100010011 : color = 12'hf63;
15'b0000101001100010100 : color = 12'he73;
15'b0000101001100010101 : color = 12'he73;
15'b0000101001100010110 : color = 12'hf30;
15'b0000101001100010111 : color = 12'hf11;
15'b0000101001100011000 : color = 12'hf73;
15'b0000101001100011001 : color = 12'he73;
15'b0000101001100011010 : color = 12'he73;
15'b0000101001100011011 : color = 12'he73;
15'b0000101001100011100 : color = 12'he61;
15'b0000101001100011101 : color = 12'hf00;
15'b0000101001100011110 : color = 12'hf53;
15'b0000101001100011111 : color = 12'he73;
15'b0000101001100100000 : color = 12'he73;
15'b0000101001100100001 : color = 12'he73;
15'b0000101001100100010 : color = 12'he73;
15'b0000101001100100011 : color = 12'he51;
15'b0000101001100100100 : color = 12'hf00;
15'b0000101001100100101 : color = 12'hf63;
15'b0000101001100100110 : color = 12'he73;
15'b0000101001100100111 : color = 12'he73;
15'b0000101001100101000 : color = 12'he73;
15'b0000101001100101001 : color = 12'he73;
15'b0000101001100101010 : color = 12'he73;
15'b0000101001100101011 : color = 12'he73;
15'b0000101001100101100 : color = 12'he73;
15'b0000101001100101101 : color = 12'he73;
15'b0000101001100101110 : color = 12'he73;
15'b0000101001100101111 : color = 12'he73;
15'b0000101001100110000 : color = 12'he73;
15'b0000101001100110001 : color = 12'he73;
15'b0000101001100110010 : color = 12'he73;
15'b0000101001100110011 : color = 12'he73;
15'b0000101001100110100 : color = 12'he73;
15'b0000101001100110101 : color = 12'he73;
15'b0000101001100110110 : color = 12'he73;
15'b0000101001100110111 : color = 12'he73;
15'b0000101001100111000 : color = 12'he73;
15'b0000101001100111001 : color = 12'he73;
15'b0000101001100111010 : color = 12'he73;
15'b0000101001100111011 : color = 12'he73;
15'b0000101001100111100 : color = 12'he73;
15'b0000101001100111101 : color = 12'he51;
15'b0000101001100111110 : color = 12'hf01;
15'b0000101001100111111 : color = 12'hf73;
15'b0000101001101000000 : color = 12'he72;
15'b0000101001101000001 : color = 12'hf10;
15'b0000101001101000010 : color = 12'hf11;
15'b0000101001101000011 : color = 12'hf73;
15'b0000101001101000100 : color = 12'he73;
15'b0000101001101000101 : color = 12'he73;
15'b0000101001101000110 : color = 12'he73;
15'b0000101001101000111 : color = 12'he73;
15'b0000101001101001000 : color = 12'he73;
15'b0000101001101001001 : color = 12'he73;
15'b0000101001101001010 : color = 12'he51;
15'b0000101001101001011 : color = 12'hf00;
15'b0000101001101001100 : color = 12'hf53;
15'b0000101001101001101 : color = 12'he73;
15'b0000101001101001110 : color = 12'he73;
15'b0000101001101001111 : color = 12'he73;
15'b0000101001101010000 : color = 12'he73;
15'b0000101001101010001 : color = 12'he73;
15'b0000101001101010010 : color = 12'he73;
15'b0000101001101010011 : color = 12'he73;
15'b0000101001101010100 : color = 12'he73;
15'b0000101001101010101 : color = 12'he73;
15'b0000101001101010110 : color = 12'he73;
15'b0000101001101010111 : color = 12'he73;
15'b0000101001101011000 : color = 12'he73;
15'b0000101001101011001 : color = 12'he73;
15'b0000101001101011010 : color = 12'he73;
15'b0000101001101011011 : color = 12'he73;
15'b0000101001101011100 : color = 12'he73;
15'b0000101001101011101 : color = 12'he73;
15'b0000101001101011110 : color = 12'he73;
15'b0000101001101011111 : color = 12'he73;
15'b0000101001101100000 : color = 12'he73;
15'b0000101001101100001 : color = 12'he73;
15'b0000101001101100010 : color = 12'he73;
15'b0000101001101100011 : color = 12'he73;
15'b0000101001101100100 : color = 12'he73;
15'b0000101001101100101 : color = 12'he73;
15'b0000101001101100110 : color = 12'he73;
15'b0000101001101100111 : color = 12'he73;
15'b0000101001101101000 : color = 12'he73;
15'b0000101001101101001 : color = 12'he73;
15'b0000101001101101010 : color = 12'he73;
15'b0000101001101101011 : color = 12'hf30;
15'b0000101001101101100 : color = 12'hf11;
15'b0000101001101101101 : color = 12'hf73;
15'b0000101001101101110 : color = 12'he73;
15'b0000101001101101111 : color = 12'he73;
15'b0000101001101110000 : color = 12'he73;
15'b0000101001101110001 : color = 12'he73;
15'b0000101001101110010 : color = 12'he73;
15'b0000101001101110011 : color = 12'he73;
15'b0000101001101110100 : color = 12'he73;
15'b0000101001101110101 : color = 12'he73;
15'b0000101001101110110 : color = 12'he73;
15'b0000101001101110111 : color = 12'he73;
15'b0000101001101111000 : color = 12'he61;
15'b0000101001101111001 : color = 12'hf52;
15'b0000101001101111010 : color = 12'he73;
15'b0000101001101111011 : color = 12'he73;
15'b0000101001101111100 : color = 12'he73;
15'b0000101001101111101 : color = 12'he73;
15'b0000101001101111110 : color = 12'he73;
15'b0000101001101111111 : color = 12'he73;
15'b0000101001110000000 : color = 12'he73;
15'b0000101001110000001 : color = 12'he73;
15'b0000101001110000010 : color = 12'he73;
15'b0000101001110000011 : color = 12'he73;
15'b0000101001110000100 : color = 12'he73;
15'b0000101001110000101 : color = 12'he73;
15'b0000101001110000110 : color = 12'he73;
15'b0000101001110000111 : color = 12'he73;
15'b0000101001110001000 : color = 12'he73;
15'b0000101001110001001 : color = 12'he73;
15'b0000101001110001010 : color = 12'he73;
15'b0000101001110001011 : color = 12'he73;
15'b0000101001110001100 : color = 12'he73;
15'b0000101001110001101 : color = 12'he73;
15'b0000101001110001110 : color = 12'he73;
15'b0000101001110001111 : color = 12'he73;
15'b0000101001110010000 : color = 12'he73;
15'b0000101001110010001 : color = 12'he73;
15'b0000101001110010010 : color = 12'he73;
15'b0000101001110010011 : color = 12'he73;
15'b0000101001110010100 : color = 12'he73;
15'b0000101001110010101 : color = 12'he72;
15'b0000101001110010110 : color = 12'hf10;
15'b0000101001110010111 : color = 12'hf32;
15'b0000101001110011000 : color = 12'he62;
15'b0000101001110011001 : color = 12'hf41;
15'b0000101001110011010 : color = 12'hf11;
15'b0000101001110011011 : color = 12'hf52;
15'b0000101001110011100 : color = 12'hf51;
15'b0000101001110011101 : color = 12'hf31;
15'b0000101001110011110 : color = 12'hf31;
15'b0000101001110011111 : color = 12'hf31;
15'b0000101001110100000 : color = 12'hf31;
15'b0000101001110100001 : color = 12'hf31;
15'b0000101001110100010 : color = 12'hf10;
15'b0000101001110100011 : color = 12'hf10;
15'b0000101001110100100 : color = 12'hf31;
15'b0000101001110100101 : color = 12'hf31;
15'b0000101001110100110 : color = 12'hf31;
15'b0000101001110100111 : color = 12'hf00;
15'b0000101001110101000 : color = 12'hf00;
15'b0000101001110101001 : color = 12'hf11;
15'b0000101001110101010 : color = 12'hf73;
15'b0000101001110101011 : color = 12'he73;
15'b0000101001110101100 : color = 12'he73;
15'b0000101001110101101 : color = 12'he73;
15'b0000101001110101110 : color = 12'he73;
15'b0000101001110101111 : color = 12'he73;
15'b0000101001110110000 : color = 12'he73;
15'b0000101001110110001 : color = 12'he73;
15'b0000101001110110010 : color = 12'he73;
15'b0000101001110110011 : color = 12'he73;
15'b0000101001110110100 : color = 12'he73;
15'b0000101001110110101 : color = 12'he73;
15'b0000101001110110110 : color = 12'he73;
15'b0000101001110110111 : color = 12'he73;
15'b0000101001110111000 : color = 12'he73;
15'b0000101001110111001 : color = 12'he73;
15'b0000101001110111010 : color = 12'he73;
15'b0000101001110111011 : color = 12'he73;
15'b0000101001110111100 : color = 12'he73;
15'b0000101001110111101 : color = 12'he73;
15'b0000101001110111110 : color = 12'he73;
15'b0000101001110111111 : color = 12'he73;
15'b0000101001111000000 : color = 12'he73;
15'b0000101001111000001 : color = 12'he73;
15'b0000101001111000010 : color = 12'he73;
15'b0000101001111000011 : color = 12'he73;
15'b0000101001111000100 : color = 12'he61;
15'b0000101001111000101 : color = 12'hf00;
15'b0000101001111000110 : color = 12'hf00;
15'b0000101001111000111 : color = 12'hf11;
15'b0000101001111001000 : color = 12'hf73;
15'b0000101001111001001 : color = 12'he73;
15'b0000101001111001010 : color = 12'he51;
15'b0000101001111001011 : color = 12'hf00;
15'b0000101001111001100 : color = 12'hf53;
15'b0000101001111001101 : color = 12'he73;
15'b0000101001111001110 : color = 12'he73;
15'b0000101001111001111 : color = 12'hf40;
15'b0000101001111010000 : color = 12'hf00;
15'b0000101001111010001 : color = 12'hf42;
15'b0000101001111010010 : color = 12'hf73;
15'b0000101001111010011 : color = 12'he73;
15'b0000101001111010100 : color = 12'he73;
15'b0000101001111010101 : color = 12'he73;
15'b0000101001111010110 : color = 12'he73;
15'b0000101001111010111 : color = 12'he73;
15'b0000101001111011000 : color = 12'he73;
15'b0000101001111011001 : color = 12'he73;
15'b0000101001111011010 : color = 12'he73;
15'b0000101001111011011 : color = 12'he73;
15'b0000101001111011100 : color = 12'he73;
15'b0000101001111011101 : color = 12'he73;
15'b0000101001111011110 : color = 12'he73;
15'b0000101001111011111 : color = 12'he73;
15'b0000101001111100000 : color = 12'he73;
15'b0000101001111100001 : color = 12'he73;
15'b0000101001111100010 : color = 12'he73;
15'b0000101001111100011 : color = 12'he73;
15'b0000101001111100100 : color = 12'he73;
15'b0000101001111100101 : color = 12'he73;
15'b0000101001111100110 : color = 12'he73;
15'b0000101001111100111 : color = 12'he73;
15'b0000101001111101000 : color = 12'he73;
15'b0000101001111101001 : color = 12'he73;
15'b0000101001111101010 : color = 12'he73;
15'b0000101001111101011 : color = 12'he73;
15'b0000101001111101100 : color = 12'he73;
15'b0000101001111101101 : color = 12'he73;
15'b0000101001111101110 : color = 12'he73;
15'b0000101001111101111 : color = 12'he73;
15'b0000101001111110000 : color = 12'he73;
15'b0000101001111110001 : color = 12'hf62;
15'b0000101001111110010 : color = 12'hf31;
15'b0000101001111110011 : color = 12'hf11;
15'b0000101001111110100 : color = 12'hf63;
15'b0000101001111110101 : color = 12'he73;
15'b0000101001111110110 : color = 12'he73;
15'b0000101001111110111 : color = 12'hf40;
15'b0000101001111111000 : color = 12'hf01;
15'b0000101001111111001 : color = 12'hf73;
15'b0000101001111111010 : color = 12'he73;
15'b0000101001111111011 : color = 12'he73;
15'b0000101001111111100 : color = 12'hf30;
15'b0000101001111111101 : color = 12'hf11;
15'b0000101001111111110 : color = 12'hf73;
15'b0000101001111111111 : color = 12'he73;
15'b0000101010000000000 : color = 12'he73;
15'b0000101010000000001 : color = 12'he73;
15'b0000101010000000010 : color = 12'he73;
15'b0000101010000000011 : color = 12'he73;
15'b0000101010000000100 : color = 12'he73;
15'b0000101010000000101 : color = 12'he73;
15'b0000101010000000110 : color = 12'he73;
15'b0000101010000000111 : color = 12'he73;
15'b0000101010000001000 : color = 12'he73;
15'b0000101010000001001 : color = 12'he73;
15'b0000101010000001010 : color = 12'he73;
15'b0000101010000001011 : color = 12'he73;
15'b0000101010000001100 : color = 12'he73;
15'b0000101010000001101 : color = 12'he73;
15'b0000101010000001110 : color = 12'he73;
15'b0000101010000001111 : color = 12'he73;
15'b0000101010000010000 : color = 12'he73;
15'b0000101010000010001 : color = 12'he73;
15'b0000101010000010010 : color = 12'he73;
15'b0000101010000010011 : color = 12'he73;
15'b0000101001001010010 : color = 12'he73;
15'b0000101001001010011 : color = 12'he73;
15'b0000101001001010100 : color = 12'he73;
15'b0000101001001010101 : color = 12'he73;
15'b0000101001001010110 : color = 12'he73;
15'b0000101001001010111 : color = 12'he73;
15'b0000101001001011000 : color = 12'he73;
15'b0000101001001011001 : color = 12'he73;
15'b0000101001001011010 : color = 12'he73;
15'b0000101001001011011 : color = 12'he73;
15'b0000101001001011100 : color = 12'he51;
15'b0000101001001011101 : color = 12'hf11;
15'b0000101001001011110 : color = 12'hf73;
15'b0000101001001011111 : color = 12'he73;
15'b0000101001001100000 : color = 12'he73;
15'b0000101001001100001 : color = 12'he73;
15'b0000101001001100010 : color = 12'he73;
15'b0000101001001100011 : color = 12'he51;
15'b0000101001001100100 : color = 12'hf00;
15'b0000101001001100101 : color = 12'hf53;
15'b0000101001001100110 : color = 12'he73;
15'b0000101001001100111 : color = 12'he61;
15'b0000101001001101000 : color = 12'hf00;
15'b0000101001001101001 : color = 12'hf42;
15'b0000101001001101010 : color = 12'he73;
15'b0000101001001101011 : color = 12'he73;
15'b0000101001001101100 : color = 12'he73;
15'b0000101001001101101 : color = 12'he73;
15'b0000101001001101110 : color = 12'hf40;
15'b0000101001001101111 : color = 12'hf00;
15'b0000101001001110000 : color = 12'hf63;
15'b0000101001001110001 : color = 12'he73;
15'b0000101001001110010 : color = 12'he73;
15'b0000101001001110011 : color = 12'he73;
15'b0000101001001110100 : color = 12'he73;
15'b0000101001001110101 : color = 12'he73;
15'b0000101001001110110 : color = 12'he73;
15'b0000101001001110111 : color = 12'he73;
15'b0000101001001111000 : color = 12'he73;
15'b0000101001001111001 : color = 12'he73;
15'b0000101001001111010 : color = 12'he73;
15'b0000101001001111011 : color = 12'he73;
15'b0000101001001111100 : color = 12'he73;
15'b0000101001001111101 : color = 12'he73;
15'b0000101001001111110 : color = 12'he73;
15'b0000101001001111111 : color = 12'he73;
15'b0000101001010000000 : color = 12'he73;
15'b0000101001010000001 : color = 12'he73;
15'b0000101001010000010 : color = 12'he73;
15'b0000101001010000011 : color = 12'he73;
15'b0000101001010000100 : color = 12'he73;
15'b0000101001010000101 : color = 12'he73;
15'b0000101001010000110 : color = 12'he73;
15'b0000101001010000111 : color = 12'he73;
15'b0000101001010001000 : color = 12'he62;
15'b0000101001010001001 : color = 12'hf10;
15'b0000101001010001010 : color = 12'hf11;
15'b0000101001010001011 : color = 12'hf41;
15'b0000101001010001100 : color = 12'hf11;
15'b0000101001010001101 : color = 12'hf63;
15'b0000101001010001110 : color = 12'he73;
15'b0000101001010001111 : color = 12'he73;
15'b0000101001010010000 : color = 12'he73;
15'b0000101001010010001 : color = 12'he73;
15'b0000101001010010010 : color = 12'he73;
15'b0000101001010010011 : color = 12'he73;
15'b0000101001010010100 : color = 12'he73;
15'b0000101001010010101 : color = 12'he73;
15'b0000101001010010110 : color = 12'he72;
15'b0000101001010010111 : color = 12'hf00;
15'b0000101001010011000 : color = 12'hf32;
15'b0000101001010011001 : color = 12'he73;
15'b0000101001010011010 : color = 12'he73;
15'b0000101001010011011 : color = 12'he73;
15'b0000101001010011100 : color = 12'he73;
15'b0000101001010011101 : color = 12'he73;
15'b0000101001010011110 : color = 12'he73;
15'b0000101001010011111 : color = 12'he73;
15'b0000101001010100000 : color = 12'he73;
15'b0000101001010100001 : color = 12'he73;
15'b0000101001010100010 : color = 12'he73;
15'b0000101001010100011 : color = 12'he73;
15'b0000101001010100100 : color = 12'he73;
15'b0000101001010100101 : color = 12'he73;
15'b0000101001010100110 : color = 12'he73;
15'b0000101001010100111 : color = 12'he73;
15'b0000101001010101000 : color = 12'he73;
15'b0000101001010101001 : color = 12'he73;
15'b0000101001010101010 : color = 12'he73;
15'b0000101001010101011 : color = 12'he73;
15'b0000101001010101100 : color = 12'he73;
15'b0000101001010101101 : color = 12'he73;
15'b0000101001010101110 : color = 12'he73;
15'b0000101001010101111 : color = 12'he73;
15'b0000101001010110000 : color = 12'he73;
15'b0000101001010110001 : color = 12'he73;
15'b0000101001010110010 : color = 12'he73;
15'b0000101001010110011 : color = 12'he73;
15'b0000101001010110100 : color = 12'he73;
15'b0000101001010110101 : color = 12'he73;
15'b0000101001010110110 : color = 12'he73;
15'b0000101001010110111 : color = 12'he73;
15'b0000101001010111000 : color = 12'he61;
15'b0000101001010111001 : color = 12'hf00;
15'b0000101001010111010 : color = 12'hf42;
15'b0000101001010111011 : color = 12'he73;
15'b0000101001010111100 : color = 12'he73;
15'b0000101001010111101 : color = 12'he73;
15'b0000101001010111110 : color = 12'hf40;
15'b0000101001010111111 : color = 12'hf00;
15'b0000101001011000000 : color = 12'hf53;
15'b0000101001011000001 : color = 12'he73;
15'b0000101001011000010 : color = 12'he73;
15'b0000101001011000011 : color = 12'he73;
15'b0000101001011000100 : color = 12'he61;
15'b0000101001011000101 : color = 12'hf00;
15'b0000101001011000110 : color = 12'hf00;
15'b0000101001011000111 : color = 12'hf52;
15'b0000101001011001000 : color = 12'he73;
15'b0000101001011001001 : color = 12'he73;
15'b0000101001011001010 : color = 12'he73;
15'b0000101001011001011 : color = 12'he73;
15'b0000101001011001100 : color = 12'he73;
15'b0000101001011001101 : color = 12'he73;
15'b0000101001011001110 : color = 12'he73;
15'b0000101001011001111 : color = 12'he73;
15'b0000101001011010000 : color = 12'he73;
15'b0000101001011010001 : color = 12'he73;
15'b0000101001011010010 : color = 12'he73;
15'b0000101001011010011 : color = 12'he73;
15'b0000101001011010100 : color = 12'he73;
15'b0000101001011010101 : color = 12'he73;
15'b0000101001011010110 : color = 12'he73;
15'b0000101001011010111 : color = 12'he73;
15'b0000101001011011000 : color = 12'he73;
15'b0000101001011011001 : color = 12'he73;
15'b0000101001011011010 : color = 12'he73;
15'b0000101001011011011 : color = 12'he73;
15'b0000101001011011100 : color = 12'he73;
15'b0000101001011011101 : color = 12'he73;
15'b0000101001011011110 : color = 12'he73;
15'b0000101001011011111 : color = 12'he73;
15'b0000101001011100000 : color = 12'he73;
15'b0000101001011100001 : color = 12'he73;
15'b0000101001011100010 : color = 12'he73;
15'b0000101001011100011 : color = 12'he73;
15'b0000101001011100100 : color = 12'he73;
15'b0000101001011100101 : color = 12'he72;
15'b0000101001011100110 : color = 12'hf00;
15'b0000101001011100111 : color = 12'hf42;
15'b0000101001011101000 : color = 12'he73;
15'b0000101001011101001 : color = 12'he73;
15'b0000101001011101010 : color = 12'he73;
15'b0000101001011101011 : color = 12'he73;
15'b0000101001011101100 : color = 12'he73;
15'b0000101001011101101 : color = 12'he73;
15'b0000101001011101110 : color = 12'he73;
15'b0000101001011101111 : color = 12'he72;
15'b0000101001011110000 : color = 12'hf32;
15'b0000101001011110001 : color = 12'hf63;
15'b0000101001011110010 : color = 12'he73;
15'b0000101001011110011 : color = 12'he73;
15'b0000101001011110100 : color = 12'he73;
15'b0000101001011110101 : color = 12'hf40;
15'b0000101001011110110 : color = 12'hf01;
15'b0000101001011110111 : color = 12'hf73;
15'b0000101001011111000 : color = 12'he73;
15'b0000101001011111001 : color = 12'he73;
15'b0000101001011111010 : color = 12'he73;
15'b0000101001011111011 : color = 12'he73;
15'b0000101001011111100 : color = 12'he73;
15'b0000101001011111101 : color = 12'he73;
15'b0000101001011111110 : color = 12'he73;
15'b0000101001011111111 : color = 12'he73;
15'b0000101001100000000 : color = 12'he73;
15'b0000101001100000001 : color = 12'he73;
15'b0000101001100000010 : color = 12'he73;
15'b0000101001100000011 : color = 12'he73;
15'b0000101001100000100 : color = 12'he73;
15'b0000101001100000101 : color = 12'he73;
15'b0000101001100000110 : color = 12'he73;
15'b0000101001100000111 : color = 12'he73;
15'b0000101001100001000 : color = 12'he73;
15'b0000101001100001001 : color = 12'he73;
15'b0000101001100001010 : color = 12'he73;
15'b0000101001100001011 : color = 12'he73;
15'b0000101001100001100 : color = 12'he73;
15'b0000101001100001101 : color = 12'he73;
15'b0000101001100001110 : color = 12'he73;
15'b0000101001100001111 : color = 12'he73;
15'b0000101001100010000 : color = 12'he73;
15'b0000101001100010001 : color = 12'he73;
15'b0000101001100010010 : color = 12'he73;
15'b0000101001100010011 : color = 12'he73;
15'b0000101001100010100 : color = 12'he73;
15'b0000101001100010101 : color = 12'he72;
15'b0000101001100010110 : color = 12'hf10;
15'b0000101001100010111 : color = 12'hf00;
15'b0000101001100011000 : color = 12'hf53;
15'b0000101001100011001 : color = 12'he73;
15'b0000101001100011010 : color = 12'he73;
15'b0000101001100011011 : color = 12'he73;
15'b0000101001100011100 : color = 12'he73;
15'b0000101001100011101 : color = 12'he73;
15'b0000101001100011110 : color = 12'he73;
15'b0000101001100011111 : color = 12'he73;
15'b0000101001100100000 : color = 12'he73;
15'b0000101001100100001 : color = 12'he73;
15'b0000101001100100010 : color = 12'he73;
15'b0000101001100100011 : color = 12'he73;
15'b0000101001100100100 : color = 12'he73;
15'b0000101001100100101 : color = 12'he73;
15'b0000101001100100110 : color = 12'he73;
15'b0000101001100100111 : color = 12'he73;
15'b0000101001100101000 : color = 12'he73;
15'b0000101001100101001 : color = 12'he73;
15'b0000101001100101010 : color = 12'he73;
15'b0000101001100101011 : color = 12'he73;
15'b0000101001100101100 : color = 12'he73;
15'b0000101001100101101 : color = 12'he73;
15'b0000101001100101110 : color = 12'he73;
15'b0000101001100101111 : color = 12'he73;
15'b0000101001100110000 : color = 12'he73;
15'b0000101001100110001 : color = 12'he73;
15'b0000101001100110010 : color = 12'he73;
15'b0000101001100110011 : color = 12'he73;
15'b0000101001100110100 : color = 12'he73;
15'b0000101001100110101 : color = 12'he73;
15'b0000101001100110110 : color = 12'he73;
15'b0000101001100110111 : color = 12'he73;
15'b0000101001100111000 : color = 12'he73;
15'b0000101001100111001 : color = 12'he73;
15'b0000101001100111010 : color = 12'he51;
15'b0000101001100111011 : color = 12'hf00;
15'b0000101001100111100 : color = 12'hf63;
15'b0000101001100111101 : color = 12'he73;
15'b0000101001100111110 : color = 12'he73;
15'b0000101001100111111 : color = 12'hf30;
15'b0000101001101000000 : color = 12'hf11;
15'b0000101001101000001 : color = 12'hf73;
15'b0000101001101000010 : color = 12'he73;
15'b0000101001101000011 : color = 12'he73;
15'b0000101001101000100 : color = 12'he73;
15'b0000101001101000101 : color = 12'he61;
15'b0000101001101000110 : color = 12'hf00;
15'b0000101001101000111 : color = 12'hf53;
15'b0000101001101001000 : color = 12'he72;
15'b0000101001101001001 : color = 12'hf41;
15'b0000101001101001010 : color = 12'hf31;
15'b0000101001101001011 : color = 12'hf31;
15'b0000101001101001100 : color = 12'hf10;
15'b0000101001101001101 : color = 12'hf00;
15'b0000101001101001110 : color = 12'hf63;
15'b0000101001101001111 : color = 12'he73;
15'b0000101001101010000 : color = 12'he73;
15'b0000101001101010001 : color = 12'he73;
15'b0000101001101010010 : color = 12'he73;
15'b0000101001101010011 : color = 12'he73;
15'b0000101001101010100 : color = 12'he73;
15'b0000101001101010101 : color = 12'he73;
15'b0000101001101010110 : color = 12'he73;
15'b0000101001101010111 : color = 12'he73;
15'b0000101001101011000 : color = 12'he73;
15'b0000101001101011001 : color = 12'he73;
15'b0000101001101011010 : color = 12'he73;
15'b0000101001101011011 : color = 12'he73;
15'b0000101001101011100 : color = 12'he73;
15'b0000101001101011101 : color = 12'he73;
15'b0000101001101011110 : color = 12'he73;
15'b0000101001101011111 : color = 12'he73;
15'b0000101001101100000 : color = 12'he73;
15'b0000101001101100001 : color = 12'he73;
15'b0000101001101100010 : color = 12'he73;
15'b0000101001101100011 : color = 12'he73;
15'b0000101001101100100 : color = 12'he73;
15'b0000101001101100101 : color = 12'he73;
15'b0000101001101100110 : color = 12'hf30;
15'b0000101001101100111 : color = 12'hf32;
15'b0000101001101101000 : color = 12'he73;
15'b0000101001101101001 : color = 12'he73;
15'b0000101001101101010 : color = 12'he61;
15'b0000101001101101011 : color = 12'hf00;
15'b0000101001101101100 : color = 12'hf32;
15'b0000101001101101101 : color = 12'he73;
15'b0000101001101101110 : color = 12'he73;
15'b0000101001101101111 : color = 12'he73;
15'b0000101001101110000 : color = 12'he73;
15'b0000101001101110001 : color = 12'he73;
15'b0000101001101110010 : color = 12'he73;
15'b0000101001101110011 : color = 12'he51;
15'b0000101001101110100 : color = 12'hf00;
15'b0000101001101110101 : color = 12'hf53;
15'b0000101001101110110 : color = 12'he73;
15'b0000101001101110111 : color = 12'he73;
15'b0000101001101111000 : color = 12'he73;
15'b0000101001101111001 : color = 12'he73;
15'b0000101001101111010 : color = 12'he73;
15'b0000101001101111011 : color = 12'he73;
15'b0000101001101111100 : color = 12'he73;
15'b0000101001101111101 : color = 12'he73;
15'b0000101001101111110 : color = 12'he73;
15'b0000101001101111111 : color = 12'he73;
15'b0000101001110000000 : color = 12'he73;
15'b0000101001110000001 : color = 12'he73;
15'b0000101001110000010 : color = 12'he73;
15'b0000101001110000011 : color = 12'he73;
15'b0000101001110000100 : color = 12'he73;
15'b0000101001110000101 : color = 12'he73;
15'b0000101001110000110 : color = 12'he73;
15'b0000101001110000111 : color = 12'he73;
15'b0000101001110001000 : color = 12'he73;
15'b0000101001110001001 : color = 12'he73;
15'b0000101001110001010 : color = 12'he73;
15'b0000101001110001011 : color = 12'he73;
15'b0000101001110001100 : color = 12'he73;
15'b0000101001110001101 : color = 12'he73;
15'b0000101001110001110 : color = 12'he73;
15'b0000101001110001111 : color = 12'he73;
15'b0000101001110010000 : color = 12'he73;
15'b0000101001110010001 : color = 12'he73;
15'b0000101001110010010 : color = 12'he73;
15'b0000101001110010011 : color = 12'he73;
15'b0000101001110010100 : color = 12'hf30;
15'b0000101001110010101 : color = 12'hf00;
15'b0000101001110010110 : color = 12'hf31;
15'b0000101001110010111 : color = 12'hf31;
15'b0000101001110011000 : color = 12'hf31;
15'b0000101001110011001 : color = 12'hf31;
15'b0000101001110011010 : color = 12'hf31;
15'b0000101001110011011 : color = 12'hf31;
15'b0000101001110011100 : color = 12'hf31;
15'b0000101001110011101 : color = 12'hf31;
15'b0000101001110011110 : color = 12'hf31;
15'b0000101001110011111 : color = 12'hf31;
15'b0000101001110100000 : color = 12'hf31;
15'b0000101001110100001 : color = 12'hf00;
15'b0000101001110100010 : color = 12'hf00;
15'b0000101001110100011 : color = 12'hf53;
15'b0000101001110100100 : color = 12'he73;
15'b0000101001110100101 : color = 12'he73;
15'b0000101001110100110 : color = 12'he73;
15'b0000101001110100111 : color = 12'he73;
15'b0000101001110101000 : color = 12'he73;
15'b0000101001110101001 : color = 12'he73;
15'b0000101001110101010 : color = 12'he73;
15'b0000101001110101011 : color = 12'he73;
15'b0000101001110101100 : color = 12'he73;
15'b0000101001110101101 : color = 12'he73;
15'b0000101001110101110 : color = 12'he73;
15'b0000101001110101111 : color = 12'he73;
15'b0000101001110110000 : color = 12'he73;
15'b0000101001110110001 : color = 12'he73;
15'b0000101001110110010 : color = 12'he73;
15'b0000101001110110011 : color = 12'he73;
15'b0000101001110110100 : color = 12'he73;
15'b0000101001110110101 : color = 12'he73;
15'b0000101001110110110 : color = 12'he73;
15'b0000101001110110111 : color = 12'he73;
15'b0000101001110111000 : color = 12'he73;
15'b0000101001110111001 : color = 12'he73;
15'b0000101001110111010 : color = 12'he73;
15'b0000101001110111011 : color = 12'he73;
15'b0000101001110111100 : color = 12'he73;
15'b0000101001110111101 : color = 12'he73;
15'b0000101001110111110 : color = 12'he62;
15'b0000101001110111111 : color = 12'hf10;
15'b0000101001111000000 : color = 12'hf00;
15'b0000101001111000001 : color = 12'hf11;
15'b0000101001111000010 : color = 12'hf52;
15'b0000101001111000011 : color = 12'he73;
15'b0000101001111000100 : color = 12'he73;
15'b0000101001111000101 : color = 12'he72;
15'b0000101001111000110 : color = 12'hf62;
15'b0000101001111000111 : color = 12'he73;
15'b0000101001111001000 : color = 12'he73;
15'b0000101001111001001 : color = 12'he73;
15'b0000101001111001010 : color = 12'he73;
15'b0000101001111001011 : color = 12'hf30;
15'b0000101001111001100 : color = 12'hf32;
15'b0000101001111001101 : color = 12'he73;
15'b0000101001111001110 : color = 12'he73;
15'b0000101001111001111 : color = 12'he73;
15'b0000101001111010000 : color = 12'he73;
15'b0000101001111010001 : color = 12'he73;
15'b0000101001111010010 : color = 12'he73;
15'b0000101001111010011 : color = 12'he73;
15'b0000101001111010100 : color = 12'he73;
15'b0000101001111010101 : color = 12'he73;
15'b0000101001111010110 : color = 12'he73;
15'b0000101001111010111 : color = 12'he73;
15'b0000101001111011000 : color = 12'he73;
15'b0000101001111011001 : color = 12'he73;
15'b0000101001111011010 : color = 12'he73;
15'b0000101001111011011 : color = 12'he73;
15'b0000101001111011100 : color = 12'he73;
15'b0000101001111011101 : color = 12'he73;
15'b0000101001111011110 : color = 12'he73;
15'b0000101001111011111 : color = 12'he73;
15'b0000101001111100000 : color = 12'he73;
15'b0000101001111100001 : color = 12'he73;
15'b0000101001111100010 : color = 12'he73;
15'b0000101001111100011 : color = 12'he73;
15'b0000101001111100100 : color = 12'he73;
15'b0000101001111100101 : color = 12'he73;
15'b0000101001111100110 : color = 12'he73;
15'b0000101001111100111 : color = 12'he73;
15'b0000101001111101000 : color = 12'he73;
15'b0000101001111101001 : color = 12'he73;
15'b0000101001111101010 : color = 12'he73;
15'b0000101001111101011 : color = 12'he73;
15'b0000101001111101100 : color = 12'he72;
15'b0000101001111101101 : color = 12'hf00;
15'b0000101001111101110 : color = 12'hf00;
15'b0000101001111101111 : color = 12'hf52;
15'b0000101001111110000 : color = 12'he73;
15'b0000101001111110001 : color = 12'he73;
15'b0000101001111110010 : color = 12'he73;
15'b0000101001111110011 : color = 12'he51;
15'b0000101001111110100 : color = 12'hf00;
15'b0000101001111110101 : color = 12'hf53;
15'b0000101001111110110 : color = 12'he73;
15'b0000101001111110111 : color = 12'he73;
15'b0000101001111111000 : color = 12'he73;
15'b0000101001111111001 : color = 12'hf51;
15'b0000101001111111010 : color = 12'hf00;
15'b0000101001111111011 : color = 12'hf00;
15'b0000101001111111100 : color = 12'hf52;
15'b0000101001111111101 : color = 12'hf73;
15'b0000101001111111110 : color = 12'he73;
15'b0000101001111111111 : color = 12'he73;
15'b0000101010000000000 : color = 12'he73;
15'b0000101010000000001 : color = 12'he73;
15'b0000101010000000010 : color = 12'he73;
15'b0000101010000000011 : color = 12'he73;
15'b0000101010000000100 : color = 12'he73;
15'b0000101010000000101 : color = 12'he73;
15'b0000101010000000110 : color = 12'he73;
15'b0000101010000000111 : color = 12'he73;
15'b0000101010000001000 : color = 12'he73;
15'b0000101010000001001 : color = 12'he73;
15'b0000101010000001010 : color = 12'he73;
15'b0000101010000001011 : color = 12'he73;
15'b0000101010000001100 : color = 12'he73;
15'b0000101010000001101 : color = 12'he73;
15'b0000101010000001110 : color = 12'he73;
15'b0000101010000001111 : color = 12'he73;
15'b0000101010000010000 : color = 12'he73;
15'b0000101010000010001 : color = 12'he73;
15'b0000101010000010010 : color = 12'he73;
15'b0000101010000010011 : color = 12'he73;
15'b0000101010000010100 : color = 12'he73;
15'b0000101010000010101 : color = 12'he73;
15'b0000101010000010110 : color = 12'hf62;
15'b0000101010000010111 : color = 12'hf41;
15'b0000101010000011000 : color = 12'hf10;
15'b0000101010000011001 : color = 12'hf00;
15'b0000101010000011010 : color = 12'hf32;
15'b0000101010000011011 : color = 12'hf63;
15'b0000101010000011100 : color = 12'he73;
15'b0000101010000011101 : color = 12'he73;
15'b0000101010000011110 : color = 12'he73;
15'b0000101010000011111 : color = 12'he72;
15'b0000101010000100000 : color = 12'hf10;
15'b0000101010000100001 : color = 12'hf11;
15'b0000101010000100010 : color = 12'hf73;
15'b0000101010000100011 : color = 12'he73;
15'b0000101010000100100 : color = 12'he73;
15'b0000101010000100101 : color = 12'hf30;
15'b0000101010000100110 : color = 12'hf11;
15'b0000101010000100111 : color = 12'hf73;
15'b0000101010000101000 : color = 12'he73;
15'b0000101010000101001 : color = 12'he73;
15'b0000101010000101010 : color = 12'he62;
15'b0000101010000101011 : color = 12'hf63;
15'b0000101010000101100 : color = 12'he73;
15'b0000101010000101101 : color = 12'he73;
15'b0000101010000101110 : color = 12'he73;
15'b0000101010000101111 : color = 12'he73;
15'b0000101010000110000 : color = 12'he73;
15'b0000101010000110001 : color = 12'he73;
15'b0000101010000110010 : color = 12'he73;
15'b0000101010000110011 : color = 12'he73;
15'b0000101010000110100 : color = 12'he73;
15'b0000101010000110101 : color = 12'he73;
15'b0000101010000110110 : color = 12'he73;
15'b0000101010000110111 : color = 12'he73;
15'b0000101010000111000 : color = 12'he73;
15'b0000101010000111001 : color = 12'he73;
15'b0000101010000111010 : color = 12'he73;
15'b0000101010000111011 : color = 12'he73;
15'b0000101010000111100 : color = 12'he73;
15'b0000101001001111011 : color = 12'he73;
15'b0000101001001111100 : color = 12'he73;
15'b0000101001001111101 : color = 12'he73;
15'b0000101001001111110 : color = 12'he73;
15'b0000101001001111111 : color = 12'he73;
15'b0000101001010000000 : color = 12'he73;
15'b0000101001010000001 : color = 12'he73;
15'b0000101001010000010 : color = 12'he73;
15'b0000101001010000011 : color = 12'he73;
15'b0000101001010000100 : color = 12'he61;
15'b0000101001010000101 : color = 12'hf11;
15'b0000101001010000110 : color = 12'hf73;
15'b0000101001010000111 : color = 12'he73;
15'b0000101001010001000 : color = 12'he73;
15'b0000101001010001001 : color = 12'he73;
15'b0000101001010001010 : color = 12'he73;
15'b0000101001010001011 : color = 12'he73;
15'b0000101001010001100 : color = 12'he72;
15'b0000101001010001101 : color = 12'hf31;
15'b0000101001010001110 : color = 12'hf73;
15'b0000101001010001111 : color = 12'he72;
15'b0000101001010010000 : color = 12'hf10;
15'b0000101001010010001 : color = 12'hf32;
15'b0000101001010010010 : color = 12'he73;
15'b0000101001010010011 : color = 12'he73;
15'b0000101001010010100 : color = 12'he73;
15'b0000101001010010101 : color = 12'he73;
15'b0000101001010010110 : color = 12'he73;
15'b0000101001010010111 : color = 12'he72;
15'b0000101001010011000 : color = 12'hf00;
15'b0000101001010011001 : color = 12'hf01;
15'b0000101001010011010 : color = 12'hf73;
15'b0000101001010011011 : color = 12'he73;
15'b0000101001010011100 : color = 12'he73;
15'b0000101001010011101 : color = 12'he73;
15'b0000101001010011110 : color = 12'he73;
15'b0000101001010011111 : color = 12'he73;
15'b0000101001010100000 : color = 12'he73;
15'b0000101001010100001 : color = 12'he73;
15'b0000101001010100010 : color = 12'he73;
15'b0000101001010100011 : color = 12'he73;
15'b0000101001010100100 : color = 12'he73;
15'b0000101001010100101 : color = 12'he73;
15'b0000101001010100110 : color = 12'he73;
15'b0000101001010100111 : color = 12'he73;
15'b0000101001010101000 : color = 12'he73;
15'b0000101001010101001 : color = 12'he73;
15'b0000101001010101010 : color = 12'he73;
15'b0000101001010101011 : color = 12'he73;
15'b0000101001010101100 : color = 12'he73;
15'b0000101001010101101 : color = 12'he73;
15'b0000101001010101110 : color = 12'he73;
15'b0000101001010101111 : color = 12'he72;
15'b0000101001010110000 : color = 12'hf30;
15'b0000101001010110001 : color = 12'hf00;
15'b0000101001010110010 : color = 12'hf32;
15'b0000101001010110011 : color = 12'hf73;
15'b0000101001010110100 : color = 12'he73;
15'b0000101001010110101 : color = 12'he62;
15'b0000101001010110110 : color = 12'hf10;
15'b0000101001010110111 : color = 12'hf52;
15'b0000101001010111000 : color = 12'he73;
15'b0000101001010111001 : color = 12'he73;
15'b0000101001010111010 : color = 12'he73;
15'b0000101001010111011 : color = 12'he73;
15'b0000101001010111100 : color = 12'he73;
15'b0000101001010111101 : color = 12'he73;
15'b0000101001010111110 : color = 12'he73;
15'b0000101001010111111 : color = 12'he72;
15'b0000101001011000000 : color = 12'hf00;
15'b0000101001011000001 : color = 12'hf32;
15'b0000101001011000010 : color = 12'he73;
15'b0000101001011000011 : color = 12'he73;
15'b0000101001011000100 : color = 12'he73;
15'b0000101001011000101 : color = 12'he73;
15'b0000101001011000110 : color = 12'he73;
15'b0000101001011000111 : color = 12'he73;
15'b0000101001011001000 : color = 12'he73;
15'b0000101001011001001 : color = 12'he73;
15'b0000101001011001010 : color = 12'he73;
15'b0000101001011001011 : color = 12'he73;
15'b0000101001011001100 : color = 12'he73;
15'b0000101001011001101 : color = 12'he73;
15'b0000101001011001110 : color = 12'he73;
15'b0000101001011001111 : color = 12'he73;
15'b0000101001011010000 : color = 12'he73;
15'b0000101001011010001 : color = 12'he73;
15'b0000101001011010010 : color = 12'he73;
15'b0000101001011010011 : color = 12'he73;
15'b0000101001011010100 : color = 12'he73;
15'b0000101001011010101 : color = 12'he73;
15'b0000101001011010110 : color = 12'he73;
15'b0000101001011010111 : color = 12'he73;
15'b0000101001011011000 : color = 12'he73;
15'b0000101001011011001 : color = 12'he73;
15'b0000101001011011010 : color = 12'he73;
15'b0000101001011011011 : color = 12'he73;
15'b0000101001011011100 : color = 12'he73;
15'b0000101001011011101 : color = 12'he73;
15'b0000101001011011110 : color = 12'he73;
15'b0000101001011011111 : color = 12'he73;
15'b0000101001011100000 : color = 12'he61;
15'b0000101001011100001 : color = 12'hf00;
15'b0000101001011100010 : color = 12'hf42;
15'b0000101001011100011 : color = 12'he73;
15'b0000101001011100100 : color = 12'he73;
15'b0000101001011100101 : color = 12'he73;
15'b0000101001011100110 : color = 12'he73;
15'b0000101001011100111 : color = 12'hf40;
15'b0000101001011101000 : color = 12'hf00;
15'b0000101001011101001 : color = 12'hf53;
15'b0000101001011101010 : color = 12'he73;
15'b0000101001011101011 : color = 12'he73;
15'b0000101001011101100 : color = 12'he73;
15'b0000101001011101101 : color = 12'he73;
15'b0000101001011101110 : color = 12'he51;
15'b0000101001011101111 : color = 12'hf00;
15'b0000101001011110000 : color = 12'hf00;
15'b0000101001011110001 : color = 12'hf31;
15'b0000101001011110010 : color = 12'hf63;
15'b0000101001011110011 : color = 12'he73;
15'b0000101001011110100 : color = 12'he73;
15'b0000101001011110101 : color = 12'he73;
15'b0000101001011110110 : color = 12'he73;
15'b0000101001011110111 : color = 12'he73;
15'b0000101001011111000 : color = 12'he73;
15'b0000101001011111001 : color = 12'he73;
15'b0000101001011111010 : color = 12'he73;
15'b0000101001011111011 : color = 12'he73;
15'b0000101001011111100 : color = 12'he73;
15'b0000101001011111101 : color = 12'he73;
15'b0000101001011111110 : color = 12'he73;
15'b0000101001011111111 : color = 12'he73;
15'b0000101001100000000 : color = 12'he73;
15'b0000101001100000001 : color = 12'he73;
15'b0000101001100000010 : color = 12'he73;
15'b0000101001100000011 : color = 12'he73;
15'b0000101001100000100 : color = 12'he73;
15'b0000101001100000101 : color = 12'he73;
15'b0000101001100000110 : color = 12'he73;
15'b0000101001100000111 : color = 12'he73;
15'b0000101001100001000 : color = 12'he73;
15'b0000101001100001001 : color = 12'he73;
15'b0000101001100001010 : color = 12'he73;
15'b0000101001100001011 : color = 12'he73;
15'b0000101001100001100 : color = 12'he73;
15'b0000101001100001101 : color = 12'he73;
15'b0000101001100001110 : color = 12'he72;
15'b0000101001100001111 : color = 12'hf00;
15'b0000101001100010000 : color = 12'hf42;
15'b0000101001100010001 : color = 12'he73;
15'b0000101001100010010 : color = 12'he73;
15'b0000101001100010011 : color = 12'he72;
15'b0000101001100010100 : color = 12'hf52;
15'b0000101001100010101 : color = 12'hf41;
15'b0000101001100010110 : color = 12'hf31;
15'b0000101001100010111 : color = 12'hf73;
15'b0000101001100011000 : color = 12'he73;
15'b0000101001100011001 : color = 12'he73;
15'b0000101001100011010 : color = 12'he73;
15'b0000101001100011011 : color = 12'he73;
15'b0000101001100011100 : color = 12'he73;
15'b0000101001100011101 : color = 12'he73;
15'b0000101001100011110 : color = 12'hf40;
15'b0000101001100011111 : color = 12'hf01;
15'b0000101001100100000 : color = 12'hf73;
15'b0000101001100100001 : color = 12'he73;
15'b0000101001100100010 : color = 12'he73;
15'b0000101001100100011 : color = 12'he73;
15'b0000101001100100100 : color = 12'he73;
15'b0000101001100100101 : color = 12'he73;
15'b0000101001100100110 : color = 12'he73;
15'b0000101001100100111 : color = 12'he73;
15'b0000101001100101000 : color = 12'he73;
15'b0000101001100101001 : color = 12'he73;
15'b0000101001100101010 : color = 12'he73;
15'b0000101001100101011 : color = 12'he73;
15'b0000101001100101100 : color = 12'he73;
15'b0000101001100101101 : color = 12'he73;
15'b0000101001100101110 : color = 12'he73;
15'b0000101001100101111 : color = 12'he73;
15'b0000101001100110000 : color = 12'he73;
15'b0000101001100110001 : color = 12'he73;
15'b0000101001100110010 : color = 12'he73;
15'b0000101001100110011 : color = 12'he73;
15'b0000101001100110100 : color = 12'he73;
15'b0000101001100110101 : color = 12'he73;
15'b0000101001100110110 : color = 12'he73;
15'b0000101001100110111 : color = 12'he73;
15'b0000101001100111000 : color = 12'he73;
15'b0000101001100111001 : color = 12'he73;
15'b0000101001100111010 : color = 12'he73;
15'b0000101001100111011 : color = 12'he73;
15'b0000101001100111100 : color = 12'he73;
15'b0000101001100111101 : color = 12'he62;
15'b0000101001100111110 : color = 12'hf10;
15'b0000101001100111111 : color = 12'hf11;
15'b0000101001101000000 : color = 12'hf30;
15'b0000101001101000001 : color = 12'hf00;
15'b0000101001101000010 : color = 12'hf42;
15'b0000101001101000011 : color = 12'hf73;
15'b0000101001101000100 : color = 12'he73;
15'b0000101001101000101 : color = 12'he73;
15'b0000101001101000110 : color = 12'he73;
15'b0000101001101000111 : color = 12'he73;
15'b0000101001101001000 : color = 12'he73;
15'b0000101001101001001 : color = 12'he73;
15'b0000101001101001010 : color = 12'he73;
15'b0000101001101001011 : color = 12'he73;
15'b0000101001101001100 : color = 12'he73;
15'b0000101001101001101 : color = 12'he73;
15'b0000101001101001110 : color = 12'he73;
15'b0000101001101001111 : color = 12'he73;
15'b0000101001101010000 : color = 12'he73;
15'b0000101001101010001 : color = 12'he73;
15'b0000101001101010010 : color = 12'he73;
15'b0000101001101010011 : color = 12'he73;
15'b0000101001101010100 : color = 12'he73;
15'b0000101001101010101 : color = 12'he73;
15'b0000101001101010110 : color = 12'he73;
15'b0000101001101010111 : color = 12'he73;
15'b0000101001101011000 : color = 12'he73;
15'b0000101001101011001 : color = 12'he73;
15'b0000101001101011010 : color = 12'he73;
15'b0000101001101011011 : color = 12'he73;
15'b0000101001101011100 : color = 12'he73;
15'b0000101001101011101 : color = 12'he73;
15'b0000101001101011110 : color = 12'he73;
15'b0000101001101011111 : color = 12'he73;
15'b0000101001101100000 : color = 12'he73;
15'b0000101001101100001 : color = 12'he62;
15'b0000101001101100010 : color = 12'hf10;
15'b0000101001101100011 : color = 12'hf11;
15'b0000101001101100100 : color = 12'hf51;
15'b0000101001101100101 : color = 12'hf11;
15'b0000101001101100110 : color = 12'hf63;
15'b0000101001101100111 : color = 12'he73;
15'b0000101001101101000 : color = 12'hf30;
15'b0000101001101101001 : color = 12'hf42;
15'b0000101001101101010 : color = 12'he73;
15'b0000101001101101011 : color = 12'he73;
15'b0000101001101101100 : color = 12'he73;
15'b0000101001101101101 : color = 12'he73;
15'b0000101001101101110 : color = 12'he62;
15'b0000101001101101111 : color = 12'hf42;
15'b0000101001101110000 : color = 12'hf73;
15'b0000101001101110001 : color = 12'he73;
15'b0000101001101110010 : color = 12'he73;
15'b0000101001101110011 : color = 12'he62;
15'b0000101001101110100 : color = 12'hf10;
15'b0000101001101110101 : color = 12'hf00;
15'b0000101001101110110 : color = 12'hf11;
15'b0000101001101110111 : color = 12'hf73;
15'b0000101001101111000 : color = 12'he73;
15'b0000101001101111001 : color = 12'he73;
15'b0000101001101111010 : color = 12'he73;
15'b0000101001101111011 : color = 12'he73;
15'b0000101001101111100 : color = 12'he73;
15'b0000101001101111101 : color = 12'he73;
15'b0000101001101111110 : color = 12'he73;
15'b0000101001101111111 : color = 12'he73;
15'b0000101001110000000 : color = 12'he73;
15'b0000101001110000001 : color = 12'he73;
15'b0000101001110000010 : color = 12'he73;
15'b0000101001110000011 : color = 12'he73;
15'b0000101001110000100 : color = 12'he73;
15'b0000101001110000101 : color = 12'he73;
15'b0000101001110000110 : color = 12'he73;
15'b0000101001110000111 : color = 12'he73;
15'b0000101001110001000 : color = 12'he73;
15'b0000101001110001001 : color = 12'he73;
15'b0000101001110001010 : color = 12'he73;
15'b0000101001110001011 : color = 12'he73;
15'b0000101001110001100 : color = 12'he73;
15'b0000101001110001101 : color = 12'he73;
15'b0000101001110001110 : color = 12'he61;
15'b0000101001110001111 : color = 12'hf00;
15'b0000101001110010000 : color = 12'hf63;
15'b0000101001110010001 : color = 12'he73;
15'b0000101001110010010 : color = 12'he73;
15'b0000101001110010011 : color = 12'he73;
15'b0000101001110010100 : color = 12'hf30;
15'b0000101001110010101 : color = 12'hf01;
15'b0000101001110010110 : color = 12'hf73;
15'b0000101001110010111 : color = 12'he73;
15'b0000101001110011000 : color = 12'he73;
15'b0000101001110011001 : color = 12'he73;
15'b0000101001110011010 : color = 12'he73;
15'b0000101001110011011 : color = 12'he73;
15'b0000101001110011100 : color = 12'he51;
15'b0000101001110011101 : color = 12'hf00;
15'b0000101001110011110 : color = 12'hf53;
15'b0000101001110011111 : color = 12'he73;
15'b0000101001110100000 : color = 12'he73;
15'b0000101001110100001 : color = 12'he73;
15'b0000101001110100010 : color = 12'he73;
15'b0000101001110100011 : color = 12'he73;
15'b0000101001110100100 : color = 12'he73;
15'b0000101001110100101 : color = 12'he73;
15'b0000101001110100110 : color = 12'he73;
15'b0000101001110100111 : color = 12'he73;
15'b0000101001110101000 : color = 12'he73;
15'b0000101001110101001 : color = 12'he73;
15'b0000101001110101010 : color = 12'he73;
15'b0000101001110101011 : color = 12'he73;
15'b0000101001110101100 : color = 12'he73;
15'b0000101001110101101 : color = 12'he73;
15'b0000101001110101110 : color = 12'he73;
15'b0000101001110101111 : color = 12'he73;
15'b0000101001110110000 : color = 12'he73;
15'b0000101001110110001 : color = 12'he73;
15'b0000101001110110010 : color = 12'he73;
15'b0000101001110110011 : color = 12'he73;
15'b0000101001110110100 : color = 12'he73;
15'b0000101001110110101 : color = 12'he73;
15'b0000101001110110110 : color = 12'he73;
15'b0000101001110110111 : color = 12'he73;
15'b0000101001110111000 : color = 12'he73;
15'b0000101001110111001 : color = 12'he73;
15'b0000101001110111010 : color = 12'he73;
15'b0000101001110111011 : color = 12'he73;
15'b0000101001110111100 : color = 12'he73;
15'b0000101001110111101 : color = 12'hf30;
15'b0000101001110111110 : color = 12'hf11;
15'b0000101001110111111 : color = 12'hf73;
15'b0000101001111000000 : color = 12'he73;
15'b0000101001111000001 : color = 12'he73;
15'b0000101001111000010 : color = 12'he73;
15'b0000101001111000011 : color = 12'he73;
15'b0000101001111000100 : color = 12'he73;
15'b0000101001111000101 : color = 12'he73;
15'b0000101001111000110 : color = 12'he73;
15'b0000101001111000111 : color = 12'he73;
15'b0000101001111001000 : color = 12'he73;
15'b0000101001111001001 : color = 12'he72;
15'b0000101001111001010 : color = 12'hf10;
15'b0000101001111001011 : color = 12'hf32;
15'b0000101001111001100 : color = 12'he73;
15'b0000101001111001101 : color = 12'he73;
15'b0000101001111001110 : color = 12'he73;
15'b0000101001111001111 : color = 12'he73;
15'b0000101001111010000 : color = 12'he73;
15'b0000101001111010001 : color = 12'he73;
15'b0000101001111010010 : color = 12'he73;
15'b0000101001111010011 : color = 12'he73;
15'b0000101001111010100 : color = 12'he73;
15'b0000101001111010101 : color = 12'he73;
15'b0000101001111010110 : color = 12'he73;
15'b0000101001111010111 : color = 12'he73;
15'b0000101001111011000 : color = 12'he73;
15'b0000101001111011001 : color = 12'he73;
15'b0000101001111011010 : color = 12'he73;
15'b0000101001111011011 : color = 12'he73;
15'b0000101001111011100 : color = 12'he73;
15'b0000101001111011101 : color = 12'he73;
15'b0000101001111011110 : color = 12'he73;
15'b0000101001111011111 : color = 12'he73;
15'b0000101001111100000 : color = 12'he73;
15'b0000101001111100001 : color = 12'he73;
15'b0000101001111100010 : color = 12'he73;
15'b0000101001111100011 : color = 12'he73;
15'b0000101001111100100 : color = 12'hf52;
15'b0000101001111100101 : color = 12'hf30;
15'b0000101001111100110 : color = 12'hf00;
15'b0000101001111100111 : color = 12'hf00;
15'b0000101001111101000 : color = 12'hf11;
15'b0000101001111101001 : color = 12'hf63;
15'b0000101001111101010 : color = 12'he73;
15'b0000101001111101011 : color = 12'he73;
15'b0000101001111101100 : color = 12'he73;
15'b0000101001111101101 : color = 12'he73;
15'b0000101001111101110 : color = 12'he73;
15'b0000101001111101111 : color = 12'he73;
15'b0000101001111110000 : color = 12'he73;
15'b0000101001111110001 : color = 12'he73;
15'b0000101001111110010 : color = 12'he73;
15'b0000101001111110011 : color = 12'he73;
15'b0000101001111110100 : color = 12'hf30;
15'b0000101001111110101 : color = 12'hf32;
15'b0000101001111110110 : color = 12'he73;
15'b0000101001111110111 : color = 12'he73;
15'b0000101001111111000 : color = 12'he73;
15'b0000101001111111001 : color = 12'he73;
15'b0000101001111111010 : color = 12'he73;
15'b0000101001111111011 : color = 12'he73;
15'b0000101001111111100 : color = 12'he73;
15'b0000101001111111101 : color = 12'he73;
15'b0000101001111111110 : color = 12'he73;
15'b0000101001111111111 : color = 12'he73;
15'b0000101010000000000 : color = 12'he73;
15'b0000101010000000001 : color = 12'he73;
15'b0000101010000000010 : color = 12'he73;
15'b0000101010000000011 : color = 12'he73;
15'b0000101010000000100 : color = 12'he73;
15'b0000101010000000101 : color = 12'he73;
15'b0000101010000000110 : color = 12'he73;
15'b0000101010000000111 : color = 12'he73;
15'b0000101010000001000 : color = 12'he73;
15'b0000101010000001001 : color = 12'he73;
15'b0000101010000001010 : color = 12'he73;
15'b0000101010000001011 : color = 12'he73;
15'b0000101010000001100 : color = 12'he73;
15'b0000101010000001101 : color = 12'he73;
15'b0000101010000001110 : color = 12'he73;
15'b0000101010000001111 : color = 12'he73;
15'b0000101010000010000 : color = 12'he73;
15'b0000101010000010001 : color = 12'he73;
15'b0000101010000010010 : color = 12'he73;
15'b0000101010000010011 : color = 12'he73;
15'b0000101010000010100 : color = 12'he72;
15'b0000101010000010101 : color = 12'hf10;
15'b0000101010000010110 : color = 12'hf11;
15'b0000101010000010111 : color = 12'hf63;
15'b0000101010000011000 : color = 12'he73;
15'b0000101010000011001 : color = 12'he73;
15'b0000101010000011010 : color = 12'he73;
15'b0000101010000011011 : color = 12'he73;
15'b0000101010000011100 : color = 12'he51;
15'b0000101010000011101 : color = 12'hf00;
15'b0000101010000011110 : color = 12'hf53;
15'b0000101010000011111 : color = 12'he73;
15'b0000101010000100000 : color = 12'he73;
15'b0000101010000100001 : color = 12'he73;
15'b0000101010000100010 : color = 12'he73;
15'b0000101010000100011 : color = 12'he51;
15'b0000101010000100100 : color = 12'hf00;
15'b0000101010000100101 : color = 12'hf00;
15'b0000101010000100110 : color = 12'hf11;
15'b0000101010000100111 : color = 12'hf73;
15'b0000101010000101000 : color = 12'he73;
15'b0000101010000101001 : color = 12'he73;
15'b0000101010000101010 : color = 12'he73;
15'b0000101010000101011 : color = 12'he73;
15'b0000101010000101100 : color = 12'he73;
15'b0000101010000101101 : color = 12'he73;
15'b0000101010000101110 : color = 12'he73;
15'b0000101010000101111 : color = 12'he73;
15'b0000101010000110000 : color = 12'he73;
15'b0000101010000110001 : color = 12'he73;
15'b0000101010000110010 : color = 12'he73;
15'b0000101010000110011 : color = 12'he73;
15'b0000101010000110100 : color = 12'he73;
15'b0000101010000110101 : color = 12'he73;
15'b0000101010000110110 : color = 12'he73;
15'b0000101010000110111 : color = 12'he73;
15'b0000101010000111000 : color = 12'he73;
15'b0000101010000111001 : color = 12'he73;
15'b0000101010000111010 : color = 12'he73;
15'b0000101010000111011 : color = 12'he72;
15'b0000101010000111100 : color = 12'hf30;
15'b0000101010000111101 : color = 12'hf10;
15'b0000101010000111110 : color = 12'hf00;
15'b0000101010000111111 : color = 12'hf00;
15'b0000101010001000000 : color = 12'hf10;
15'b0000101010001000001 : color = 12'hf52;
15'b0000101010001000010 : color = 12'hf73;
15'b0000101010001000011 : color = 12'he73;
15'b0000101010001000100 : color = 12'he73;
15'b0000101010001000101 : color = 12'he73;
15'b0000101010001000110 : color = 12'he73;
15'b0000101010001000111 : color = 12'he73;
15'b0000101010001001000 : color = 12'he61;
15'b0000101010001001001 : color = 12'hf00;
15'b0000101010001001010 : color = 12'hf42;
15'b0000101010001001011 : color = 12'he73;
15'b0000101010001001100 : color = 12'he73;
15'b0000101010001001101 : color = 12'he73;
15'b0000101010001001110 : color = 12'hf30;
15'b0000101010001001111 : color = 12'hf11;
15'b0000101010001010000 : color = 12'hf73;
15'b0000101010001010001 : color = 12'he73;
15'b0000101010001010010 : color = 12'he73;
15'b0000101010001010011 : color = 12'he61;
15'b0000101010001010100 : color = 12'hf42;
15'b0000101010001010101 : color = 12'he73;
15'b0000101010001010110 : color = 12'he73;
15'b0000101010001010111 : color = 12'he73;
15'b0000101010001011000 : color = 12'he73;
15'b0000101010001011001 : color = 12'he73;
15'b0000101010001011010 : color = 12'he73;
15'b0000101010001011011 : color = 12'he73;
15'b0000101010001011100 : color = 12'he73;
15'b0000101010001011101 : color = 12'he73;
15'b0000101010001011110 : color = 12'he73;
15'b0000101010001011111 : color = 12'he73;
15'b0000101010001100000 : color = 12'he73;
15'b0000101010001100001 : color = 12'he73;
15'b0000101010001100010 : color = 12'he73;
15'b0000101010001100011 : color = 12'he73;
15'b0000101010001100100 : color = 12'he73;
15'b0000101010001100101 : color = 12'he73;
15'b0000101001010100100 : color = 12'he73;
15'b0000101001010100101 : color = 12'he73;
15'b0000101001010100110 : color = 12'he73;
15'b0000101001010100111 : color = 12'he73;
15'b0000101001010101000 : color = 12'he73;
15'b0000101001010101001 : color = 12'he73;
15'b0000101001010101010 : color = 12'he73;
15'b0000101001010101011 : color = 12'he73;
15'b0000101001010101100 : color = 12'he72;
15'b0000101001010101101 : color = 12'hf11;
15'b0000101001010101110 : color = 12'hf73;
15'b0000101001010101111 : color = 12'he73;
15'b0000101001010110000 : color = 12'he73;
15'b0000101001010110001 : color = 12'he73;
15'b0000101001010110010 : color = 12'he73;
15'b0000101001010110011 : color = 12'he73;
15'b0000101001010110100 : color = 12'he73;
15'b0000101001010110101 : color = 12'he73;
15'b0000101001010110110 : color = 12'he73;
15'b0000101001010110111 : color = 12'he72;
15'b0000101001010111000 : color = 12'hf10;
15'b0000101001010111001 : color = 12'hf32;
15'b0000101001010111010 : color = 12'hf73;
15'b0000101001010111011 : color = 12'he73;
15'b0000101001010111100 : color = 12'he73;
15'b0000101001010111101 : color = 12'he73;
15'b0000101001010111110 : color = 12'he73;
15'b0000101001010111111 : color = 12'he73;
15'b0000101001011000000 : color = 12'he73;
15'b0000101001011000001 : color = 12'he51;
15'b0000101001011000010 : color = 12'hf00;
15'b0000101001011000011 : color = 12'hf11;
15'b0000101001011000100 : color = 12'hf63;
15'b0000101001011000101 : color = 12'he73;
15'b0000101001011000110 : color = 12'he73;
15'b0000101001011000111 : color = 12'he73;
15'b0000101001011001000 : color = 12'he73;
15'b0000101001011001001 : color = 12'he73;
15'b0000101001011001010 : color = 12'he73;
15'b0000101001011001011 : color = 12'he73;
15'b0000101001011001100 : color = 12'he73;
15'b0000101001011001101 : color = 12'he73;
15'b0000101001011001110 : color = 12'he73;
15'b0000101001011001111 : color = 12'he73;
15'b0000101001011010000 : color = 12'he73;
15'b0000101001011010001 : color = 12'he73;
15'b0000101001011010010 : color = 12'he73;
15'b0000101001011010011 : color = 12'he73;
15'b0000101001011010100 : color = 12'he73;
15'b0000101001011010101 : color = 12'he73;
15'b0000101001011010110 : color = 12'he73;
15'b0000101001011010111 : color = 12'he72;
15'b0000101001011011000 : color = 12'hf30;
15'b0000101001011011001 : color = 12'hf00;
15'b0000101001011011010 : color = 12'hf32;
15'b0000101001011011011 : color = 12'hf73;
15'b0000101001011011100 : color = 12'he73;
15'b0000101001011011101 : color = 12'he73;
15'b0000101001011011110 : color = 12'he73;
15'b0000101001011011111 : color = 12'he62;
15'b0000101001011100000 : color = 12'hf10;
15'b0000101001011100001 : color = 12'hf10;
15'b0000101001011100010 : color = 12'hf42;
15'b0000101001011100011 : color = 12'hf62;
15'b0000101001011100100 : color = 12'he73;
15'b0000101001011100101 : color = 12'he73;
15'b0000101001011100110 : color = 12'he73;
15'b0000101001011100111 : color = 12'he73;
15'b0000101001011101000 : color = 12'he72;
15'b0000101001011101001 : color = 12'hf00;
15'b0000101001011101010 : color = 12'hf52;
15'b0000101001011101011 : color = 12'he73;
15'b0000101001011101100 : color = 12'he73;
15'b0000101001011101101 : color = 12'he73;
15'b0000101001011101110 : color = 12'he73;
15'b0000101001011101111 : color = 12'he73;
15'b0000101001011110000 : color = 12'he73;
15'b0000101001011110001 : color = 12'he73;
15'b0000101001011110010 : color = 12'hf63;
15'b0000101001011110011 : color = 12'he73;
15'b0000101001011110100 : color = 12'he73;
15'b0000101001011110101 : color = 12'he73;
15'b0000101001011110110 : color = 12'he73;
15'b0000101001011110111 : color = 12'he73;
15'b0000101001011111000 : color = 12'he73;
15'b0000101001011111001 : color = 12'he73;
15'b0000101001011111010 : color = 12'he73;
15'b0000101001011111011 : color = 12'he73;
15'b0000101001011111100 : color = 12'he73;
15'b0000101001011111101 : color = 12'he73;
15'b0000101001011111110 : color = 12'he73;
15'b0000101001011111111 : color = 12'he73;
15'b0000101001100000000 : color = 12'he73;
15'b0000101001100000001 : color = 12'he73;
15'b0000101001100000010 : color = 12'he73;
15'b0000101001100000011 : color = 12'he73;
15'b0000101001100000100 : color = 12'he73;
15'b0000101001100000101 : color = 12'he73;
15'b0000101001100000110 : color = 12'he73;
15'b0000101001100000111 : color = 12'he73;
15'b0000101001100001000 : color = 12'hf51;
15'b0000101001100001001 : color = 12'hf00;
15'b0000101001100001010 : color = 12'hf52;
15'b0000101001100001011 : color = 12'he73;
15'b0000101001100001100 : color = 12'he73;
15'b0000101001100001101 : color = 12'he73;
15'b0000101001100001110 : color = 12'he73;
15'b0000101001100001111 : color = 12'he73;
15'b0000101001100010000 : color = 12'hf40;
15'b0000101001100010001 : color = 12'hf00;
15'b0000101001100010010 : color = 12'hf53;
15'b0000101001100010011 : color = 12'he73;
15'b0000101001100010100 : color = 12'he73;
15'b0000101001100010101 : color = 12'he73;
15'b0000101001100010110 : color = 12'he73;
15'b0000101001100010111 : color = 12'he73;
15'b0000101001100011000 : color = 12'he61;
15'b0000101001100011001 : color = 12'hf00;
15'b0000101001100011010 : color = 12'hf00;
15'b0000101001100011011 : color = 12'hf00;
15'b0000101001100011100 : color = 12'hf11;
15'b0000101001100011101 : color = 12'hf52;
15'b0000101001100011110 : color = 12'hf73;
15'b0000101001100011111 : color = 12'he73;
15'b0000101001100100000 : color = 12'he73;
15'b0000101001100100001 : color = 12'he73;
15'b0000101001100100010 : color = 12'he73;
15'b0000101001100100011 : color = 12'he73;
15'b0000101001100100100 : color = 12'he73;
15'b0000101001100100101 : color = 12'he73;
15'b0000101001100100110 : color = 12'he73;
15'b0000101001100100111 : color = 12'he73;
15'b0000101001100101000 : color = 12'he73;
15'b0000101001100101001 : color = 12'he73;
15'b0000101001100101010 : color = 12'he73;
15'b0000101001100101011 : color = 12'he73;
15'b0000101001100101100 : color = 12'he73;
15'b0000101001100101101 : color = 12'he73;
15'b0000101001100101110 : color = 12'he73;
15'b0000101001100101111 : color = 12'he73;
15'b0000101001100110000 : color = 12'he73;
15'b0000101001100110001 : color = 12'he73;
15'b0000101001100110010 : color = 12'he73;
15'b0000101001100110011 : color = 12'he73;
15'b0000101001100110100 : color = 12'he73;
15'b0000101001100110101 : color = 12'he73;
15'b0000101001100110110 : color = 12'he73;
15'b0000101001100110111 : color = 12'he62;
15'b0000101001100111000 : color = 12'hf00;
15'b0000101001100111001 : color = 12'hf11;
15'b0000101001100111010 : color = 12'hf10;
15'b0000101001100111011 : color = 12'hf00;
15'b0000101001100111100 : color = 12'hf11;
15'b0000101001100111101 : color = 12'hf42;
15'b0000101001100111110 : color = 12'hf63;
15'b0000101001100111111 : color = 12'he73;
15'b0000101001101000000 : color = 12'he73;
15'b0000101001101000001 : color = 12'he73;
15'b0000101001101000010 : color = 12'he73;
15'b0000101001101000011 : color = 12'he73;
15'b0000101001101000100 : color = 12'he73;
15'b0000101001101000101 : color = 12'he73;
15'b0000101001101000110 : color = 12'he73;
15'b0000101001101000111 : color = 12'he51;
15'b0000101001101001000 : color = 12'hf01;
15'b0000101001101001001 : color = 12'hf73;
15'b0000101001101001010 : color = 12'he73;
15'b0000101001101001011 : color = 12'he73;
15'b0000101001101001100 : color = 12'he73;
15'b0000101001101001101 : color = 12'he73;
15'b0000101001101001110 : color = 12'he73;
15'b0000101001101001111 : color = 12'he73;
15'b0000101001101010000 : color = 12'he73;
15'b0000101001101010001 : color = 12'he73;
15'b0000101001101010010 : color = 12'he73;
15'b0000101001101010011 : color = 12'he73;
15'b0000101001101010100 : color = 12'he73;
15'b0000101001101010101 : color = 12'he73;
15'b0000101001101010110 : color = 12'he73;
15'b0000101001101010111 : color = 12'he73;
15'b0000101001101011000 : color = 12'he73;
15'b0000101001101011001 : color = 12'he73;
15'b0000101001101011010 : color = 12'he73;
15'b0000101001101011011 : color = 12'he73;
15'b0000101001101011100 : color = 12'he73;
15'b0000101001101011101 : color = 12'he73;
15'b0000101001101011110 : color = 12'he73;
15'b0000101001101011111 : color = 12'he73;
15'b0000101001101100000 : color = 12'he73;
15'b0000101001101100001 : color = 12'he73;
15'b0000101001101100010 : color = 12'he73;
15'b0000101001101100011 : color = 12'he73;
15'b0000101001101100100 : color = 12'he73;
15'b0000101001101100101 : color = 12'hf41;
15'b0000101001101100110 : color = 12'hf00;
15'b0000101001101100111 : color = 12'hf32;
15'b0000101001101101000 : color = 12'hf73;
15'b0000101001101101001 : color = 12'he73;
15'b0000101001101101010 : color = 12'hf40;
15'b0000101001101101011 : color = 12'hf00;
15'b0000101001101101100 : color = 12'hf11;
15'b0000101001101101101 : color = 12'hf52;
15'b0000101001101101110 : color = 12'he73;
15'b0000101001101101111 : color = 12'he73;
15'b0000101001101110000 : color = 12'he73;
15'b0000101001101110001 : color = 12'he73;
15'b0000101001101110010 : color = 12'he73;
15'b0000101001101110011 : color = 12'he73;
15'b0000101001101110100 : color = 12'he73;
15'b0000101001101110101 : color = 12'he73;
15'b0000101001101110110 : color = 12'he73;
15'b0000101001101110111 : color = 12'he73;
15'b0000101001101111000 : color = 12'he73;
15'b0000101001101111001 : color = 12'he73;
15'b0000101001101111010 : color = 12'he73;
15'b0000101001101111011 : color = 12'he73;
15'b0000101001101111100 : color = 12'he73;
15'b0000101001101111101 : color = 12'he73;
15'b0000101001101111110 : color = 12'he73;
15'b0000101001101111111 : color = 12'he73;
15'b0000101001110000000 : color = 12'he73;
15'b0000101001110000001 : color = 12'he73;
15'b0000101001110000010 : color = 12'he73;
15'b0000101001110000011 : color = 12'he73;
15'b0000101001110000100 : color = 12'he73;
15'b0000101001110000101 : color = 12'he73;
15'b0000101001110000110 : color = 12'he73;
15'b0000101001110000111 : color = 12'he73;
15'b0000101001110001000 : color = 12'he73;
15'b0000101001110001001 : color = 12'hf41;
15'b0000101001110001010 : color = 12'hf00;
15'b0000101001110001011 : color = 12'hf11;
15'b0000101001110001100 : color = 12'hf73;
15'b0000101001110001101 : color = 12'he73;
15'b0000101001110001110 : color = 12'he72;
15'b0000101001110001111 : color = 12'hf10;
15'b0000101001110010000 : color = 12'hf42;
15'b0000101001110010001 : color = 12'hf73;
15'b0000101001110010010 : color = 12'he73;
15'b0000101001110010011 : color = 12'he73;
15'b0000101001110010100 : color = 12'he73;
15'b0000101001110010101 : color = 12'he73;
15'b0000101001110010110 : color = 12'he73;
15'b0000101001110010111 : color = 12'he73;
15'b0000101001110011000 : color = 12'he73;
15'b0000101001110011001 : color = 12'he73;
15'b0000101001110011010 : color = 12'he73;
15'b0000101001110011011 : color = 12'he73;
15'b0000101001110011100 : color = 12'he73;
15'b0000101001110011101 : color = 12'he72;
15'b0000101001110011110 : color = 12'hf32;
15'b0000101001110011111 : color = 12'hf73;
15'b0000101001110100000 : color = 12'he73;
15'b0000101001110100001 : color = 12'he73;
15'b0000101001110100010 : color = 12'he73;
15'b0000101001110100011 : color = 12'he73;
15'b0000101001110100100 : color = 12'he73;
15'b0000101001110100101 : color = 12'he73;
15'b0000101001110100110 : color = 12'he73;
15'b0000101001110100111 : color = 12'he73;
15'b0000101001110101000 : color = 12'he73;
15'b0000101001110101001 : color = 12'he73;
15'b0000101001110101010 : color = 12'he73;
15'b0000101001110101011 : color = 12'he73;
15'b0000101001110101100 : color = 12'he73;
15'b0000101001110101101 : color = 12'he73;
15'b0000101001110101110 : color = 12'he73;
15'b0000101001110101111 : color = 12'he73;
15'b0000101001110110000 : color = 12'he73;
15'b0000101001110110001 : color = 12'he73;
15'b0000101001110110010 : color = 12'he73;
15'b0000101001110110011 : color = 12'he73;
15'b0000101001110110100 : color = 12'he73;
15'b0000101001110110101 : color = 12'he73;
15'b0000101001110110110 : color = 12'he73;
15'b0000101001110110111 : color = 12'hf30;
15'b0000101001110111000 : color = 12'hf42;
15'b0000101001110111001 : color = 12'he73;
15'b0000101001110111010 : color = 12'he73;
15'b0000101001110111011 : color = 12'he73;
15'b0000101001110111100 : color = 12'he73;
15'b0000101001110111101 : color = 12'he61;
15'b0000101001110111110 : color = 12'hf32;
15'b0000101001110111111 : color = 12'he73;
15'b0000101001111000000 : color = 12'he73;
15'b0000101001111000001 : color = 12'he73;
15'b0000101001111000010 : color = 12'he73;
15'b0000101001111000011 : color = 12'he73;
15'b0000101001111000100 : color = 12'he73;
15'b0000101001111000101 : color = 12'he51;
15'b0000101001111000110 : color = 12'hf00;
15'b0000101001111000111 : color = 12'hf53;
15'b0000101001111001000 : color = 12'he73;
15'b0000101001111001001 : color = 12'he73;
15'b0000101001111001010 : color = 12'he73;
15'b0000101001111001011 : color = 12'he73;
15'b0000101001111001100 : color = 12'he73;
15'b0000101001111001101 : color = 12'he73;
15'b0000101001111001110 : color = 12'he73;
15'b0000101001111001111 : color = 12'he73;
15'b0000101001111010000 : color = 12'he73;
15'b0000101001111010001 : color = 12'he73;
15'b0000101001111010010 : color = 12'he73;
15'b0000101001111010011 : color = 12'he73;
15'b0000101001111010100 : color = 12'he73;
15'b0000101001111010101 : color = 12'he73;
15'b0000101001111010110 : color = 12'he73;
15'b0000101001111010111 : color = 12'he73;
15'b0000101001111011000 : color = 12'he73;
15'b0000101001111011001 : color = 12'he73;
15'b0000101001111011010 : color = 12'he73;
15'b0000101001111011011 : color = 12'he73;
15'b0000101001111011100 : color = 12'he73;
15'b0000101001111011101 : color = 12'he73;
15'b0000101001111011110 : color = 12'he73;
15'b0000101001111011111 : color = 12'he73;
15'b0000101001111100000 : color = 12'he73;
15'b0000101001111100001 : color = 12'he73;
15'b0000101001111100010 : color = 12'he73;
15'b0000101001111100011 : color = 12'he73;
15'b0000101001111100100 : color = 12'he73;
15'b0000101001111100101 : color = 12'he73;
15'b0000101001111100110 : color = 12'hf30;
15'b0000101001111100111 : color = 12'hf11;
15'b0000101001111101000 : color = 12'hf73;
15'b0000101001111101001 : color = 12'he73;
15'b0000101001111101010 : color = 12'he73;
15'b0000101001111101011 : color = 12'he73;
15'b0000101001111101100 : color = 12'he73;
15'b0000101001111101101 : color = 12'he73;
15'b0000101001111101110 : color = 12'he73;
15'b0000101001111101111 : color = 12'he73;
15'b0000101001111110000 : color = 12'he73;
15'b0000101001111110001 : color = 12'he73;
15'b0000101001111110010 : color = 12'he72;
15'b0000101001111110011 : color = 12'hf10;
15'b0000101001111110100 : color = 12'hf32;
15'b0000101001111110101 : color = 12'he73;
15'b0000101001111110110 : color = 12'he73;
15'b0000101001111110111 : color = 12'he73;
15'b0000101001111111000 : color = 12'he73;
15'b0000101001111111001 : color = 12'he73;
15'b0000101001111111010 : color = 12'he73;
15'b0000101001111111011 : color = 12'he73;
15'b0000101001111111100 : color = 12'he73;
15'b0000101001111111101 : color = 12'he73;
15'b0000101001111111110 : color = 12'he73;
15'b0000101001111111111 : color = 12'he73;
15'b0000101010000000000 : color = 12'he73;
15'b0000101010000000001 : color = 12'he73;
15'b0000101010000000010 : color = 12'he73;
15'b0000101010000000011 : color = 12'he73;
15'b0000101010000000100 : color = 12'he73;
15'b0000101010000000101 : color = 12'he73;
15'b0000101010000000110 : color = 12'he73;
15'b0000101010000000111 : color = 12'he73;
15'b0000101010000001000 : color = 12'he73;
15'b0000101010000001001 : color = 12'he73;
15'b0000101010000001010 : color = 12'he73;
15'b0000101010000001011 : color = 12'he73;
15'b0000101010000001100 : color = 12'he61;
15'b0000101010000001101 : color = 12'hf00;
15'b0000101010000001110 : color = 12'hf00;
15'b0000101010000001111 : color = 12'hf11;
15'b0000101010000010000 : color = 12'hf63;
15'b0000101010000010001 : color = 12'he73;
15'b0000101010000010010 : color = 12'he73;
15'b0000101010000010011 : color = 12'he73;
15'b0000101010000010100 : color = 12'he73;
15'b0000101010000010101 : color = 12'he73;
15'b0000101010000010110 : color = 12'he73;
15'b0000101010000010111 : color = 12'he73;
15'b0000101010000011000 : color = 12'he73;
15'b0000101010000011001 : color = 12'he73;
15'b0000101010000011010 : color = 12'he73;
15'b0000101010000011011 : color = 12'he73;
15'b0000101010000011100 : color = 12'he73;
15'b0000101010000011101 : color = 12'hf30;
15'b0000101010000011110 : color = 12'hf32;
15'b0000101010000011111 : color = 12'he73;
15'b0000101010000100000 : color = 12'he73;
15'b0000101010000100001 : color = 12'he73;
15'b0000101010000100010 : color = 12'he73;
15'b0000101010000100011 : color = 12'he73;
15'b0000101010000100100 : color = 12'he73;
15'b0000101010000100101 : color = 12'he73;
15'b0000101010000100110 : color = 12'he73;
15'b0000101010000100111 : color = 12'he73;
15'b0000101010000101000 : color = 12'he73;
15'b0000101010000101001 : color = 12'he73;
15'b0000101010000101010 : color = 12'he73;
15'b0000101010000101011 : color = 12'he73;
15'b0000101010000101100 : color = 12'he73;
15'b0000101010000101101 : color = 12'he73;
15'b0000101010000101110 : color = 12'he73;
15'b0000101010000101111 : color = 12'he73;
15'b0000101010000110000 : color = 12'he73;
15'b0000101010000110001 : color = 12'he73;
15'b0000101010000110010 : color = 12'he73;
15'b0000101010000110011 : color = 12'he73;
15'b0000101010000110100 : color = 12'he73;
15'b0000101010000110101 : color = 12'he73;
15'b0000101010000110110 : color = 12'he73;
15'b0000101010000110111 : color = 12'he73;
15'b0000101010000111000 : color = 12'he73;
15'b0000101010000111001 : color = 12'he73;
15'b0000101010000111010 : color = 12'he73;
15'b0000101010000111011 : color = 12'he73;
15'b0000101010000111100 : color = 12'he62;
15'b0000101010000111101 : color = 12'hf10;
15'b0000101010000111110 : color = 12'hf11;
15'b0000101010000111111 : color = 12'hf73;
15'b0000101010001000000 : color = 12'he73;
15'b0000101010001000001 : color = 12'he73;
15'b0000101010001000010 : color = 12'he73;
15'b0000101010001000011 : color = 12'he73;
15'b0000101010001000100 : color = 12'he73;
15'b0000101010001000101 : color = 12'he51;
15'b0000101010001000110 : color = 12'hf00;
15'b0000101010001000111 : color = 12'hf53;
15'b0000101010001001000 : color = 12'he73;
15'b0000101010001001001 : color = 12'he73;
15'b0000101010001001010 : color = 12'he73;
15'b0000101010001001011 : color = 12'he73;
15'b0000101010001001100 : color = 12'he73;
15'b0000101010001001101 : color = 12'he51;
15'b0000101010001001110 : color = 12'hf00;
15'b0000101010001001111 : color = 12'hf00;
15'b0000101010001010000 : color = 12'hf11;
15'b0000101010001010001 : color = 12'hf73;
15'b0000101010001010010 : color = 12'he73;
15'b0000101010001010011 : color = 12'he73;
15'b0000101010001010100 : color = 12'he73;
15'b0000101010001010101 : color = 12'he73;
15'b0000101010001010110 : color = 12'he73;
15'b0000101010001010111 : color = 12'he73;
15'b0000101010001011000 : color = 12'he73;
15'b0000101010001011001 : color = 12'he73;
15'b0000101010001011010 : color = 12'he73;
15'b0000101010001011011 : color = 12'he73;
15'b0000101010001011100 : color = 12'he73;
15'b0000101010001011101 : color = 12'he73;
15'b0000101010001011110 : color = 12'he73;
15'b0000101010001011111 : color = 12'he73;
15'b0000101010001100000 : color = 12'he73;
15'b0000101010001100001 : color = 12'he73;
15'b0000101010001100010 : color = 12'he73;
15'b0000101010001100011 : color = 12'he73;
15'b0000101010001100100 : color = 12'he73;
15'b0000101010001100101 : color = 12'hf30;
15'b0000101010001100110 : color = 12'hf00;
15'b0000101010001100111 : color = 12'hf11;
15'b0000101010001101000 : color = 12'hf52;
15'b0000101010001101001 : color = 12'he73;
15'b0000101010001101010 : color = 12'he73;
15'b0000101010001101011 : color = 12'he73;
15'b0000101010001101100 : color = 12'he73;
15'b0000101010001101101 : color = 12'he73;
15'b0000101010001101110 : color = 12'he73;
15'b0000101010001101111 : color = 12'he73;
15'b0000101010001110000 : color = 12'he73;
15'b0000101010001110001 : color = 12'hf30;
15'b0000101010001110010 : color = 12'hf01;
15'b0000101010001110011 : color = 12'hf73;
15'b0000101010001110100 : color = 12'he73;
15'b0000101010001110101 : color = 12'he73;
15'b0000101010001110110 : color = 12'he73;
15'b0000101010001110111 : color = 12'hf30;
15'b0000101010001111000 : color = 12'hf11;
15'b0000101010001111001 : color = 12'hf73;
15'b0000101010001111010 : color = 12'he73;
15'b0000101010001111011 : color = 12'he73;
15'b0000101010001111100 : color = 12'he51;
15'b0000101010001111101 : color = 12'hf42;
15'b0000101010001111110 : color = 12'he73;
15'b0000101010001111111 : color = 12'he73;
15'b0000101010010000000 : color = 12'he73;
15'b0000101010010000001 : color = 12'he73;
15'b0000101010010000010 : color = 12'he73;
15'b0000101010010000011 : color = 12'he73;
15'b0000101010010000100 : color = 12'he73;
15'b0000101010010000101 : color = 12'he73;
15'b0000101010010000110 : color = 12'he73;
15'b0000101010010000111 : color = 12'he73;
15'b0000101010010001000 : color = 12'he73;
15'b0000101010010001001 : color = 12'he73;
15'b0000101010010001010 : color = 12'he73;
15'b0000101010010001011 : color = 12'he73;
15'b0000101010010001100 : color = 12'he73;
15'b0000101010010001101 : color = 12'he73;
15'b0000101010010001110 : color = 12'he73;
15'b0000101001011001101 : color = 12'he73;
15'b0000101001011001110 : color = 12'he73;
15'b0000101001011001111 : color = 12'he73;
15'b0000101001011010000 : color = 12'he73;
15'b0000101001011010001 : color = 12'he73;
15'b0000101001011010010 : color = 12'he73;
15'b0000101001011010011 : color = 12'he73;
15'b0000101001011010100 : color = 12'he72;
15'b0000101001011010101 : color = 12'hf41;
15'b0000101001011010110 : color = 12'hf73;
15'b0000101001011010111 : color = 12'he73;
15'b0000101001011011000 : color = 12'he73;
15'b0000101001011011001 : color = 12'he73;
15'b0000101001011011010 : color = 12'he73;
15'b0000101001011011011 : color = 12'he73;
15'b0000101001011011100 : color = 12'he73;
15'b0000101001011011101 : color = 12'he73;
15'b0000101001011011110 : color = 12'he73;
15'b0000101001011011111 : color = 12'he62;
15'b0000101001011100000 : color = 12'hf10;
15'b0000101001011100001 : color = 12'hf42;
15'b0000101001011100010 : color = 12'he73;
15'b0000101001011100011 : color = 12'he73;
15'b0000101001011100100 : color = 12'he73;
15'b0000101001011100101 : color = 12'he73;
15'b0000101001011100110 : color = 12'he73;
15'b0000101001011100111 : color = 12'he73;
15'b0000101001011101000 : color = 12'he73;
15'b0000101001011101001 : color = 12'he73;
15'b0000101001011101010 : color = 12'he73;
15'b0000101001011101011 : color = 12'hf30;
15'b0000101001011101100 : color = 12'hf00;
15'b0000101001011101101 : color = 12'hf00;
15'b0000101001011101110 : color = 12'hf52;
15'b0000101001011101111 : color = 12'he73;
15'b0000101001011110000 : color = 12'he73;
15'b0000101001011110001 : color = 12'he73;
15'b0000101001011110010 : color = 12'he73;
15'b0000101001011110011 : color = 12'he73;
15'b0000101001011110100 : color = 12'he73;
15'b0000101001011110101 : color = 12'he73;
15'b0000101001011110110 : color = 12'he73;
15'b0000101001011110111 : color = 12'he73;
15'b0000101001011111000 : color = 12'he73;
15'b0000101001011111001 : color = 12'he73;
15'b0000101001011111010 : color = 12'he73;
15'b0000101001011111011 : color = 12'he73;
15'b0000101001011111100 : color = 12'he73;
15'b0000101001011111101 : color = 12'he73;
15'b0000101001011111110 : color = 12'he73;
15'b0000101001011111111 : color = 12'he73;
15'b0000101001100000000 : color = 12'he73;
15'b0000101001100000001 : color = 12'he72;
15'b0000101001100000010 : color = 12'hf31;
15'b0000101001100000011 : color = 12'hf73;
15'b0000101001100000100 : color = 12'he73;
15'b0000101001100000101 : color = 12'he73;
15'b0000101001100000110 : color = 12'he73;
15'b0000101001100000111 : color = 12'he73;
15'b0000101001100001000 : color = 12'he73;
15'b0000101001100001001 : color = 12'he73;
15'b0000101001100001010 : color = 12'hf51;
15'b0000101001100001011 : color = 12'hf10;
15'b0000101001100001100 : color = 12'hf00;
15'b0000101001100001101 : color = 12'hf00;
15'b0000101001100001110 : color = 12'hf00;
15'b0000101001100001111 : color = 12'hf10;
15'b0000101001100010000 : color = 12'hf10;
15'b0000101001100010001 : color = 12'hf10;
15'b0000101001100010010 : color = 12'hf10;
15'b0000101001100010011 : color = 12'hf10;
15'b0000101001100010100 : color = 12'hf10;
15'b0000101001100010101 : color = 12'hf10;
15'b0000101001100010110 : color = 12'hf10;
15'b0000101001100010111 : color = 12'hf10;
15'b0000101001100011000 : color = 12'hf00;
15'b0000101001100011001 : color = 12'hf00;
15'b0000101001100011010 : color = 12'hf11;
15'b0000101001100011011 : color = 12'hf52;
15'b0000101001100011100 : color = 12'he73;
15'b0000101001100011101 : color = 12'he73;
15'b0000101001100011110 : color = 12'he73;
15'b0000101001100011111 : color = 12'he73;
15'b0000101001100100000 : color = 12'he73;
15'b0000101001100100001 : color = 12'he73;
15'b0000101001100100010 : color = 12'he73;
15'b0000101001100100011 : color = 12'he73;
15'b0000101001100100100 : color = 12'he73;
15'b0000101001100100101 : color = 12'he73;
15'b0000101001100100110 : color = 12'he73;
15'b0000101001100100111 : color = 12'he73;
15'b0000101001100101000 : color = 12'he73;
15'b0000101001100101001 : color = 12'he73;
15'b0000101001100101010 : color = 12'he73;
15'b0000101001100101011 : color = 12'he73;
15'b0000101001100101100 : color = 12'he73;
15'b0000101001100101101 : color = 12'he73;
15'b0000101001100101110 : color = 12'he73;
15'b0000101001100101111 : color = 12'he72;
15'b0000101001100110000 : color = 12'hf40;
15'b0000101001100110001 : color = 12'hf11;
15'b0000101001100110010 : color = 12'hf63;
15'b0000101001100110011 : color = 12'he73;
15'b0000101001100110100 : color = 12'he73;
15'b0000101001100110101 : color = 12'he73;
15'b0000101001100110110 : color = 12'he73;
15'b0000101001100110111 : color = 12'he73;
15'b0000101001100111000 : color = 12'he73;
15'b0000101001100111001 : color = 12'hf40;
15'b0000101001100111010 : color = 12'hf00;
15'b0000101001100111011 : color = 12'hf53;
15'b0000101001100111100 : color = 12'he73;
15'b0000101001100111101 : color = 12'he73;
15'b0000101001100111110 : color = 12'he73;
15'b0000101001100111111 : color = 12'he73;
15'b0000101001101000000 : color = 12'he73;
15'b0000101001101000001 : color = 12'he73;
15'b0000101001101000010 : color = 12'he72;
15'b0000101001101000011 : color = 12'hf30;
15'b0000101001101000100 : color = 12'hf00;
15'b0000101001101000101 : color = 12'hf00;
15'b0000101001101000110 : color = 12'hf31;
15'b0000101001101000111 : color = 12'hf52;
15'b0000101001101001000 : color = 12'he73;
15'b0000101001101001001 : color = 12'he73;
15'b0000101001101001010 : color = 12'he73;
15'b0000101001101001011 : color = 12'he73;
15'b0000101001101001100 : color = 12'he73;
15'b0000101001101001101 : color = 12'he73;
15'b0000101001101001110 : color = 12'he73;
15'b0000101001101001111 : color = 12'he73;
15'b0000101001101010000 : color = 12'he73;
15'b0000101001101010001 : color = 12'he73;
15'b0000101001101010010 : color = 12'he73;
15'b0000101001101010011 : color = 12'he73;
15'b0000101001101010100 : color = 12'he73;
15'b0000101001101010101 : color = 12'he73;
15'b0000101001101010110 : color = 12'he73;
15'b0000101001101010111 : color = 12'he73;
15'b0000101001101011000 : color = 12'he73;
15'b0000101001101011001 : color = 12'he73;
15'b0000101001101011010 : color = 12'he62;
15'b0000101001101011011 : color = 12'hf52;
15'b0000101001101011100 : color = 12'hf31;
15'b0000101001101011101 : color = 12'hf10;
15'b0000101001101011110 : color = 12'hf10;
15'b0000101001101011111 : color = 12'hf00;
15'b0000101001101100000 : color = 12'hf00;
15'b0000101001101100001 : color = 12'hf10;
15'b0000101001101100010 : color = 12'hf42;
15'b0000101001101100011 : color = 12'hf63;
15'b0000101001101100100 : color = 12'he73;
15'b0000101001101100101 : color = 12'he73;
15'b0000101001101100110 : color = 12'he73;
15'b0000101001101100111 : color = 12'he73;
15'b0000101001101101000 : color = 12'he73;
15'b0000101001101101001 : color = 12'he73;
15'b0000101001101101010 : color = 12'he73;
15'b0000101001101101011 : color = 12'he73;
15'b0000101001101101100 : color = 12'he73;
15'b0000101001101101101 : color = 12'he73;
15'b0000101001101101110 : color = 12'he73;
15'b0000101001101101111 : color = 12'he73;
15'b0000101001101110000 : color = 12'hf40;
15'b0000101001101110001 : color = 12'hf01;
15'b0000101001101110010 : color = 12'hf73;
15'b0000101001101110011 : color = 12'he73;
15'b0000101001101110100 : color = 12'he73;
15'b0000101001101110101 : color = 12'he73;
15'b0000101001101110110 : color = 12'he73;
15'b0000101001101110111 : color = 12'he73;
15'b0000101001101111000 : color = 12'he73;
15'b0000101001101111001 : color = 12'he73;
15'b0000101001101111010 : color = 12'he73;
15'b0000101001101111011 : color = 12'he73;
15'b0000101001101111100 : color = 12'he73;
15'b0000101001101111101 : color = 12'he73;
15'b0000101001101111110 : color = 12'he73;
15'b0000101001101111111 : color = 12'he73;
15'b0000101001110000000 : color = 12'he73;
15'b0000101001110000001 : color = 12'he73;
15'b0000101001110000010 : color = 12'he73;
15'b0000101001110000011 : color = 12'he73;
15'b0000101001110000100 : color = 12'he73;
15'b0000101001110000101 : color = 12'he73;
15'b0000101001110000110 : color = 12'he73;
15'b0000101001110000111 : color = 12'he73;
15'b0000101001110001000 : color = 12'he73;
15'b0000101001110001001 : color = 12'he73;
15'b0000101001110001010 : color = 12'he73;
15'b0000101001110001011 : color = 12'he73;
15'b0000101001110001100 : color = 12'he62;
15'b0000101001110001101 : color = 12'hf10;
15'b0000101001110001110 : color = 12'hf11;
15'b0000101001110001111 : color = 12'hf52;
15'b0000101001110010000 : color = 12'he73;
15'b0000101001110010001 : color = 12'he73;
15'b0000101001110010010 : color = 12'he73;
15'b0000101001110010011 : color = 12'he73;
15'b0000101001110010100 : color = 12'hf51;
15'b0000101001110010101 : color = 12'hf10;
15'b0000101001110010110 : color = 12'hf00;
15'b0000101001110010111 : color = 12'hf00;
15'b0000101001110011000 : color = 12'hf42;
15'b0000101001110011001 : color = 12'hf63;
15'b0000101001110011010 : color = 12'he73;
15'b0000101001110011011 : color = 12'he73;
15'b0000101001110011100 : color = 12'he73;
15'b0000101001110011101 : color = 12'he73;
15'b0000101001110011110 : color = 12'he73;
15'b0000101001110011111 : color = 12'he73;
15'b0000101001110100000 : color = 12'he73;
15'b0000101001110100001 : color = 12'he73;
15'b0000101001110100010 : color = 12'he73;
15'b0000101001110100011 : color = 12'he73;
15'b0000101001110100100 : color = 12'he73;
15'b0000101001110100101 : color = 12'he73;
15'b0000101001110100110 : color = 12'he73;
15'b0000101001110100111 : color = 12'he73;
15'b0000101001110101000 : color = 12'he73;
15'b0000101001110101001 : color = 12'he73;
15'b0000101001110101010 : color = 12'he73;
15'b0000101001110101011 : color = 12'he73;
15'b0000101001110101100 : color = 12'he73;
15'b0000101001110101101 : color = 12'he73;
15'b0000101001110101110 : color = 12'he73;
15'b0000101001110101111 : color = 12'he73;
15'b0000101001110110000 : color = 12'he73;
15'b0000101001110110001 : color = 12'hf30;
15'b0000101001110110010 : color = 12'hf00;
15'b0000101001110110011 : color = 12'hf01;
15'b0000101001110110100 : color = 12'hf73;
15'b0000101001110110101 : color = 12'he73;
15'b0000101001110110110 : color = 12'he73;
15'b0000101001110110111 : color = 12'he73;
15'b0000101001110111000 : color = 12'he72;
15'b0000101001110111001 : color = 12'hf30;
15'b0000101001110111010 : color = 12'hf00;
15'b0000101001110111011 : color = 12'hf31;
15'b0000101001110111100 : color = 12'hf52;
15'b0000101001110111101 : color = 12'hf62;
15'b0000101001110111110 : color = 12'hf63;
15'b0000101001110111111 : color = 12'he73;
15'b0000101001111000000 : color = 12'he73;
15'b0000101001111000001 : color = 12'he73;
15'b0000101001111000010 : color = 12'he73;
15'b0000101001111000011 : color = 12'he73;
15'b0000101001111000100 : color = 12'he73;
15'b0000101001111000101 : color = 12'he73;
15'b0000101001111000110 : color = 12'he73;
15'b0000101001111000111 : color = 12'he72;
15'b0000101001111001000 : color = 12'hf62;
15'b0000101001111001001 : color = 12'hf62;
15'b0000101001111001010 : color = 12'hf52;
15'b0000101001111001011 : color = 12'hf52;
15'b0000101001111001100 : color = 12'he73;
15'b0000101001111001101 : color = 12'he73;
15'b0000101001111001110 : color = 12'he73;
15'b0000101001111001111 : color = 12'he73;
15'b0000101001111010000 : color = 12'he73;
15'b0000101001111010001 : color = 12'he73;
15'b0000101001111010010 : color = 12'he73;
15'b0000101001111010011 : color = 12'he73;
15'b0000101001111010100 : color = 12'he73;
15'b0000101001111010101 : color = 12'he73;
15'b0000101001111010110 : color = 12'he73;
15'b0000101001111010111 : color = 12'he73;
15'b0000101001111011000 : color = 12'he73;
15'b0000101001111011001 : color = 12'he73;
15'b0000101001111011010 : color = 12'he73;
15'b0000101001111011011 : color = 12'he73;
15'b0000101001111011100 : color = 12'he73;
15'b0000101001111011101 : color = 12'he73;
15'b0000101001111011110 : color = 12'he73;
15'b0000101001111011111 : color = 12'he51;
15'b0000101001111100000 : color = 12'hf11;
15'b0000101001111100001 : color = 12'hf73;
15'b0000101001111100010 : color = 12'he73;
15'b0000101001111100011 : color = 12'he73;
15'b0000101001111100100 : color = 12'he73;
15'b0000101001111100101 : color = 12'he73;
15'b0000101001111100110 : color = 12'he73;
15'b0000101001111100111 : color = 12'he73;
15'b0000101001111101000 : color = 12'he73;
15'b0000101001111101001 : color = 12'he73;
15'b0000101001111101010 : color = 12'he73;
15'b0000101001111101011 : color = 12'he73;
15'b0000101001111101100 : color = 12'he73;
15'b0000101001111101101 : color = 12'he73;
15'b0000101001111101110 : color = 12'he51;
15'b0000101001111101111 : color = 12'hf00;
15'b0000101001111110000 : color = 12'hf53;
15'b0000101001111110001 : color = 12'he73;
15'b0000101001111110010 : color = 12'he73;
15'b0000101001111110011 : color = 12'he73;
15'b0000101001111110100 : color = 12'he73;
15'b0000101001111110101 : color = 12'he73;
15'b0000101001111110110 : color = 12'he73;
15'b0000101001111110111 : color = 12'he73;
15'b0000101001111111000 : color = 12'he73;
15'b0000101001111111001 : color = 12'he73;
15'b0000101001111111010 : color = 12'he73;
15'b0000101001111111011 : color = 12'he73;
15'b0000101001111111100 : color = 12'he73;
15'b0000101001111111101 : color = 12'he73;
15'b0000101001111111110 : color = 12'he73;
15'b0000101001111111111 : color = 12'he73;
15'b0000101010000000000 : color = 12'he73;
15'b0000101010000000001 : color = 12'he73;
15'b0000101010000000010 : color = 12'he73;
15'b0000101010000000011 : color = 12'he73;
15'b0000101010000000100 : color = 12'he73;
15'b0000101010000000101 : color = 12'he73;
15'b0000101010000000110 : color = 12'he73;
15'b0000101010000000111 : color = 12'he73;
15'b0000101010000001000 : color = 12'he73;
15'b0000101010000001001 : color = 12'he73;
15'b0000101010000001010 : color = 12'he73;
15'b0000101010000001011 : color = 12'he73;
15'b0000101010000001100 : color = 12'he73;
15'b0000101010000001101 : color = 12'he73;
15'b0000101010000001110 : color = 12'he73;
15'b0000101010000001111 : color = 12'hf30;
15'b0000101010000010000 : color = 12'hf11;
15'b0000101010000010001 : color = 12'hf73;
15'b0000101010000010010 : color = 12'he73;
15'b0000101010000010011 : color = 12'he73;
15'b0000101010000010100 : color = 12'he73;
15'b0000101010000010101 : color = 12'he73;
15'b0000101010000010110 : color = 12'he73;
15'b0000101010000010111 : color = 12'he73;
15'b0000101010000011000 : color = 12'he73;
15'b0000101010000011001 : color = 12'he73;
15'b0000101010000011010 : color = 12'he73;
15'b0000101010000011011 : color = 12'he72;
15'b0000101010000011100 : color = 12'hf10;
15'b0000101010000011101 : color = 12'hf32;
15'b0000101010000011110 : color = 12'he73;
15'b0000101010000011111 : color = 12'he73;
15'b0000101010000100000 : color = 12'he73;
15'b0000101010000100001 : color = 12'he73;
15'b0000101010000100010 : color = 12'he73;
15'b0000101010000100011 : color = 12'he73;
15'b0000101010000100100 : color = 12'he73;
15'b0000101010000100101 : color = 12'he73;
15'b0000101010000100110 : color = 12'he73;
15'b0000101010000100111 : color = 12'he73;
15'b0000101010000101000 : color = 12'he73;
15'b0000101010000101001 : color = 12'he73;
15'b0000101010000101010 : color = 12'he73;
15'b0000101010000101011 : color = 12'he73;
15'b0000101010000101100 : color = 12'he73;
15'b0000101010000101101 : color = 12'he73;
15'b0000101010000101110 : color = 12'he73;
15'b0000101010000101111 : color = 12'he73;
15'b0000101010000110000 : color = 12'he73;
15'b0000101010000110001 : color = 12'he73;
15'b0000101010000110010 : color = 12'he73;
15'b0000101010000110011 : color = 12'he73;
15'b0000101010000110100 : color = 12'he73;
15'b0000101010000110101 : color = 12'he73;
15'b0000101010000110110 : color = 12'hf41;
15'b0000101010000110111 : color = 12'hf53;
15'b0000101010000111000 : color = 12'he73;
15'b0000101010000111001 : color = 12'he73;
15'b0000101010000111010 : color = 12'he73;
15'b0000101010000111011 : color = 12'he73;
15'b0000101010000111100 : color = 12'he73;
15'b0000101010000111101 : color = 12'he73;
15'b0000101010000111110 : color = 12'he73;
15'b0000101010000111111 : color = 12'he73;
15'b0000101010001000000 : color = 12'he73;
15'b0000101010001000001 : color = 12'he73;
15'b0000101010001000010 : color = 12'he73;
15'b0000101010001000011 : color = 12'he73;
15'b0000101010001000100 : color = 12'he73;
15'b0000101010001000101 : color = 12'he73;
15'b0000101010001000110 : color = 12'hf30;
15'b0000101010001000111 : color = 12'hf32;
15'b0000101010001001000 : color = 12'he73;
15'b0000101010001001001 : color = 12'he73;
15'b0000101010001001010 : color = 12'he73;
15'b0000101010001001011 : color = 12'he73;
15'b0000101010001001100 : color = 12'he72;
15'b0000101010001001101 : color = 12'hf30;
15'b0000101010001001110 : color = 12'hf42;
15'b0000101010001001111 : color = 12'he73;
15'b0000101010001010000 : color = 12'he73;
15'b0000101010001010001 : color = 12'he73;
15'b0000101010001010010 : color = 12'he73;
15'b0000101010001010011 : color = 12'he73;
15'b0000101010001010100 : color = 12'he73;
15'b0000101010001010101 : color = 12'he73;
15'b0000101010001010110 : color = 12'he73;
15'b0000101010001010111 : color = 12'he73;
15'b0000101010001011000 : color = 12'he73;
15'b0000101010001011001 : color = 12'he73;
15'b0000101010001011010 : color = 12'he73;
15'b0000101010001011011 : color = 12'he73;
15'b0000101010001011100 : color = 12'he73;
15'b0000101010001011101 : color = 12'he73;
15'b0000101010001011110 : color = 12'he73;
15'b0000101010001011111 : color = 12'he73;
15'b0000101010001100000 : color = 12'he73;
15'b0000101010001100001 : color = 12'he73;
15'b0000101010001100010 : color = 12'he73;
15'b0000101010001100011 : color = 12'he73;
15'b0000101010001100100 : color = 12'he61;
15'b0000101010001100101 : color = 12'hf00;
15'b0000101010001100110 : color = 12'hf42;
15'b0000101010001100111 : color = 12'he73;
15'b0000101010001101000 : color = 12'he73;
15'b0000101010001101001 : color = 12'he73;
15'b0000101010001101010 : color = 12'he73;
15'b0000101010001101011 : color = 12'he73;
15'b0000101010001101100 : color = 12'he73;
15'b0000101010001101101 : color = 12'he73;
15'b0000101010001101110 : color = 12'he51;
15'b0000101010001101111 : color = 12'hf00;
15'b0000101010001110000 : color = 12'hf53;
15'b0000101010001110001 : color = 12'he73;
15'b0000101010001110010 : color = 12'he73;
15'b0000101010001110011 : color = 12'he73;
15'b0000101010001110100 : color = 12'he73;
15'b0000101010001110101 : color = 12'he73;
15'b0000101010001110110 : color = 12'he73;
15'b0000101010001110111 : color = 12'hf40;
15'b0000101010001111000 : color = 12'hf00;
15'b0000101010001111001 : color = 12'hf00;
15'b0000101010001111010 : color = 12'hf63;
15'b0000101010001111011 : color = 12'he73;
15'b0000101010001111100 : color = 12'he73;
15'b0000101010001111101 : color = 12'he73;
15'b0000101010001111110 : color = 12'he73;
15'b0000101010001111111 : color = 12'he73;
15'b0000101010010000000 : color = 12'he73;
15'b0000101010010000001 : color = 12'he73;
15'b0000101010010000010 : color = 12'he73;
15'b0000101010010000011 : color = 12'he73;
15'b0000101010010000100 : color = 12'he73;
15'b0000101010010000101 : color = 12'he73;
15'b0000101010010000110 : color = 12'he73;
15'b0000101010010000111 : color = 12'he73;
15'b0000101010010001000 : color = 12'he73;
15'b0000101010010001001 : color = 12'he73;
15'b0000101010010001010 : color = 12'he73;
15'b0000101010010001011 : color = 12'he73;
15'b0000101010010001100 : color = 12'he73;
15'b0000101010010001101 : color = 12'he73;
15'b0000101010010001110 : color = 12'he61;
15'b0000101010010001111 : color = 12'hf32;
15'b0000101010010010000 : color = 12'hf73;
15'b0000101010010010001 : color = 12'he73;
15'b0000101010010010010 : color = 12'he73;
15'b0000101010010010011 : color = 12'he73;
15'b0000101010010010100 : color = 12'he73;
15'b0000101010010010101 : color = 12'he73;
15'b0000101010010010110 : color = 12'he73;
15'b0000101010010010111 : color = 12'he73;
15'b0000101010010011000 : color = 12'he73;
15'b0000101010010011001 : color = 12'hf40;
15'b0000101010010011010 : color = 12'hf00;
15'b0000101010010011011 : color = 12'hf53;
15'b0000101010010011100 : color = 12'he73;
15'b0000101010010011101 : color = 12'he73;
15'b0000101010010011110 : color = 12'he73;
15'b0000101010010011111 : color = 12'he73;
15'b0000101010010100000 : color = 12'hf30;
15'b0000101010010100001 : color = 12'hf32;
15'b0000101010010100010 : color = 12'he73;
15'b0000101010010100011 : color = 12'he73;
15'b0000101010010100100 : color = 12'he73;
15'b0000101010010100101 : color = 12'he51;
15'b0000101010010100110 : color = 12'hf32;
15'b0000101010010100111 : color = 12'he73;
15'b0000101010010101000 : color = 12'he73;
15'b0000101010010101001 : color = 12'he73;
15'b0000101010010101010 : color = 12'he73;
15'b0000101010010101011 : color = 12'he73;
15'b0000101010010101100 : color = 12'he73;
15'b0000101010010101101 : color = 12'he73;
15'b0000101010010101110 : color = 12'he73;
15'b0000101010010101111 : color = 12'he73;
15'b0000101010010110000 : color = 12'he73;
15'b0000101010010110001 : color = 12'he73;
15'b0000101010010110010 : color = 12'he73;
15'b0000101010010110011 : color = 12'he73;
15'b0000101010010110100 : color = 12'he73;
15'b0000101010010110101 : color = 12'he73;
15'b0000101010010110110 : color = 12'he73;
15'b0000101010010110111 : color = 12'he73;
15'b0000101001011110110 : color = 12'he73;
15'b0000101001011110111 : color = 12'he73;
15'b0000101001011111000 : color = 12'he73;
15'b0000101001011111001 : color = 12'he73;
15'b0000101001011111010 : color = 12'he73;
15'b0000101001011111011 : color = 12'he73;
15'b0000101001011111100 : color = 12'he73;
15'b0000101001011111101 : color = 12'he73;
15'b0000101001011111110 : color = 12'he73;
15'b0000101001011111111 : color = 12'he73;
15'b0000101001100000000 : color = 12'he73;
15'b0000101001100000001 : color = 12'he73;
15'b0000101001100000010 : color = 12'he73;
15'b0000101001100000011 : color = 12'he73;
15'b0000101001100000100 : color = 12'he73;
15'b0000101001100000101 : color = 12'he73;
15'b0000101001100000110 : color = 12'he72;
15'b0000101001100000111 : color = 12'hf41;
15'b0000101001100001000 : color = 12'hf11;
15'b0000101001100001001 : color = 12'hf63;
15'b0000101001100001010 : color = 12'he73;
15'b0000101001100001011 : color = 12'he73;
15'b0000101001100001100 : color = 12'he73;
15'b0000101001100001101 : color = 12'he73;
15'b0000101001100001110 : color = 12'he73;
15'b0000101001100001111 : color = 12'he73;
15'b0000101001100010000 : color = 12'he73;
15'b0000101001100010001 : color = 12'he73;
15'b0000101001100010010 : color = 12'he73;
15'b0000101001100010011 : color = 12'he73;
15'b0000101001100010100 : color = 12'he72;
15'b0000101001100010101 : color = 12'hf10;
15'b0000101001100010110 : color = 12'hf00;
15'b0000101001100010111 : color = 12'hf31;
15'b0000101001100011000 : color = 12'hf62;
15'b0000101001100011001 : color = 12'he73;
15'b0000101001100011010 : color = 12'he73;
15'b0000101001100011011 : color = 12'he73;
15'b0000101001100011100 : color = 12'he73;
15'b0000101001100011101 : color = 12'he73;
15'b0000101001100011110 : color = 12'he73;
15'b0000101001100011111 : color = 12'he73;
15'b0000101001100100000 : color = 12'he73;
15'b0000101001100100001 : color = 12'he73;
15'b0000101001100100010 : color = 12'he73;
15'b0000101001100100011 : color = 12'he73;
15'b0000101001100100100 : color = 12'he73;
15'b0000101001100100101 : color = 12'he73;
15'b0000101001100100110 : color = 12'he73;
15'b0000101001100100111 : color = 12'he73;
15'b0000101001100101000 : color = 12'he73;
15'b0000101001100101001 : color = 12'he73;
15'b0000101001100101010 : color = 12'he73;
15'b0000101001100101011 : color = 12'he73;
15'b0000101001100101100 : color = 12'he73;
15'b0000101001100101101 : color = 12'he73;
15'b0000101001100101110 : color = 12'he73;
15'b0000101001100101111 : color = 12'he73;
15'b0000101001100110000 : color = 12'he73;
15'b0000101001100110001 : color = 12'he73;
15'b0000101001100110010 : color = 12'he73;
15'b0000101001100110011 : color = 12'he73;
15'b0000101001100110100 : color = 12'he73;
15'b0000101001100110101 : color = 12'he72;
15'b0000101001100110110 : color = 12'hf52;
15'b0000101001100110111 : color = 12'hf41;
15'b0000101001100111000 : color = 12'hf30;
15'b0000101001100111001 : color = 12'hf10;
15'b0000101001100111010 : color = 12'hf10;
15'b0000101001100111011 : color = 12'hf10;
15'b0000101001100111100 : color = 12'hf00;
15'b0000101001100111101 : color = 12'hf00;
15'b0000101001100111110 : color = 12'hf00;
15'b0000101001100111111 : color = 12'hf00;
15'b0000101001101000000 : color = 12'hf00;
15'b0000101001101000001 : color = 12'hf00;
15'b0000101001101000010 : color = 12'hf11;
15'b0000101001101000011 : color = 12'hf73;
15'b0000101001101000100 : color = 12'he73;
15'b0000101001101000101 : color = 12'he73;
15'b0000101001101000110 : color = 12'he73;
15'b0000101001101000111 : color = 12'he73;
15'b0000101001101001000 : color = 12'he73;
15'b0000101001101001001 : color = 12'he73;
15'b0000101001101001010 : color = 12'he73;
15'b0000101001101001011 : color = 12'he73;
15'b0000101001101001100 : color = 12'he73;
15'b0000101001101001101 : color = 12'he73;
15'b0000101001101001110 : color = 12'he73;
15'b0000101001101001111 : color = 12'he73;
15'b0000101001101010000 : color = 12'he73;
15'b0000101001101010001 : color = 12'he73;
15'b0000101001101010010 : color = 12'he73;
15'b0000101001101010011 : color = 12'he73;
15'b0000101001101010100 : color = 12'he73;
15'b0000101001101010101 : color = 12'he73;
15'b0000101001101010110 : color = 12'he73;
15'b0000101001101010111 : color = 12'he62;
15'b0000101001101011000 : color = 12'hf10;
15'b0000101001101011001 : color = 12'hf52;
15'b0000101001101011010 : color = 12'he73;
15'b0000101001101011011 : color = 12'he73;
15'b0000101001101011100 : color = 12'he73;
15'b0000101001101011101 : color = 12'he73;
15'b0000101001101011110 : color = 12'he73;
15'b0000101001101011111 : color = 12'he73;
15'b0000101001101100000 : color = 12'he73;
15'b0000101001101100001 : color = 12'he73;
15'b0000101001101100010 : color = 12'hf40;
15'b0000101001101100011 : color = 12'hf00;
15'b0000101001101100100 : color = 12'hf53;
15'b0000101001101100101 : color = 12'he73;
15'b0000101001101100110 : color = 12'he73;
15'b0000101001101100111 : color = 12'he73;
15'b0000101001101101000 : color = 12'he73;
15'b0000101001101101001 : color = 12'he73;
15'b0000101001101101010 : color = 12'he73;
15'b0000101001101101011 : color = 12'he73;
15'b0000101001101101100 : color = 12'he73;
15'b0000101001101101101 : color = 12'hf51;
15'b0000101001101101110 : color = 12'hf53;
15'b0000101001101101111 : color = 12'he73;
15'b0000101001101110000 : color = 12'he73;
15'b0000101001101110001 : color = 12'he73;
15'b0000101001101110010 : color = 12'he73;
15'b0000101001101110011 : color = 12'he73;
15'b0000101001101110100 : color = 12'he73;
15'b0000101001101110101 : color = 12'he73;
15'b0000101001101110110 : color = 12'he73;
15'b0000101001101110111 : color = 12'he73;
15'b0000101001101111000 : color = 12'he73;
15'b0000101001101111001 : color = 12'he73;
15'b0000101001101111010 : color = 12'he73;
15'b0000101001101111011 : color = 12'he73;
15'b0000101001101111100 : color = 12'he73;
15'b0000101001101111101 : color = 12'he73;
15'b0000101001101111110 : color = 12'he73;
15'b0000101001101111111 : color = 12'he73;
15'b0000101001110000000 : color = 12'he73;
15'b0000101001110000001 : color = 12'he73;
15'b0000101001110000010 : color = 12'he73;
15'b0000101001110000011 : color = 12'hf30;
15'b0000101001110000100 : color = 12'hf00;
15'b0000101001110000101 : color = 12'hf00;
15'b0000101001110000110 : color = 12'hf00;
15'b0000101001110000111 : color = 12'hf11;
15'b0000101001110001000 : color = 12'hf52;
15'b0000101001110001001 : color = 12'hf73;
15'b0000101001110001010 : color = 12'he73;
15'b0000101001110001011 : color = 12'he73;
15'b0000101001110001100 : color = 12'he73;
15'b0000101001110001101 : color = 12'he73;
15'b0000101001110001110 : color = 12'he73;
15'b0000101001110001111 : color = 12'he73;
15'b0000101001110010000 : color = 12'he73;
15'b0000101001110010001 : color = 12'he73;
15'b0000101001110010010 : color = 12'he73;
15'b0000101001110010011 : color = 12'he73;
15'b0000101001110010100 : color = 12'he62;
15'b0000101001110010101 : color = 12'hf10;
15'b0000101001110010110 : color = 12'hf10;
15'b0000101001110010111 : color = 12'hf10;
15'b0000101001110011000 : color = 12'hf10;
15'b0000101001110011001 : color = 12'hf00;
15'b0000101001110011010 : color = 12'hf01;
15'b0000101001110011011 : color = 12'hf73;
15'b0000101001110011100 : color = 12'he73;
15'b0000101001110011101 : color = 12'he73;
15'b0000101001110011110 : color = 12'he73;
15'b0000101001110011111 : color = 12'he73;
15'b0000101001110100000 : color = 12'he73;
15'b0000101001110100001 : color = 12'he73;
15'b0000101001110100010 : color = 12'he73;
15'b0000101001110100011 : color = 12'he73;
15'b0000101001110100100 : color = 12'he73;
15'b0000101001110100101 : color = 12'he73;
15'b0000101001110100110 : color = 12'he73;
15'b0000101001110100111 : color = 12'he73;
15'b0000101001110101000 : color = 12'he73;
15'b0000101001110101001 : color = 12'he73;
15'b0000101001110101010 : color = 12'he73;
15'b0000101001110101011 : color = 12'he73;
15'b0000101001110101100 : color = 12'he73;
15'b0000101001110101101 : color = 12'he73;
15'b0000101001110101110 : color = 12'he73;
15'b0000101001110101111 : color = 12'he73;
15'b0000101001110110000 : color = 12'he73;
15'b0000101001110110001 : color = 12'he73;
15'b0000101001110110010 : color = 12'he73;
15'b0000101001110110011 : color = 12'he62;
15'b0000101001110110100 : color = 12'hf10;
15'b0000101001110110101 : color = 12'hf10;
15'b0000101001110110110 : color = 12'hf52;
15'b0000101001110110111 : color = 12'he73;
15'b0000101001110111000 : color = 12'he73;
15'b0000101001110111001 : color = 12'he73;
15'b0000101001110111010 : color = 12'he73;
15'b0000101001110111011 : color = 12'he73;
15'b0000101001110111100 : color = 12'he73;
15'b0000101001110111101 : color = 12'he73;
15'b0000101001110111110 : color = 12'he72;
15'b0000101001110111111 : color = 12'hf41;
15'b0000101001111000000 : color = 12'hf00;
15'b0000101001111000001 : color = 12'hf00;
15'b0000101001111000010 : color = 12'hf00;
15'b0000101001111000011 : color = 12'hf00;
15'b0000101001111000100 : color = 12'hf10;
15'b0000101001111000101 : color = 12'hf31;
15'b0000101001111000110 : color = 12'hf31;
15'b0000101001111000111 : color = 12'hf31;
15'b0000101001111001000 : color = 12'hf42;
15'b0000101001111001001 : color = 12'hf73;
15'b0000101001111001010 : color = 12'he73;
15'b0000101001111001011 : color = 12'he73;
15'b0000101001111001100 : color = 12'he73;
15'b0000101001111001101 : color = 12'he73;
15'b0000101001111001110 : color = 12'he73;
15'b0000101001111001111 : color = 12'he73;
15'b0000101001111010000 : color = 12'he73;
15'b0000101001111010001 : color = 12'he73;
15'b0000101001111010010 : color = 12'he73;
15'b0000101001111010011 : color = 12'he73;
15'b0000101001111010100 : color = 12'he73;
15'b0000101001111010101 : color = 12'he73;
15'b0000101001111010110 : color = 12'he73;
15'b0000101001111010111 : color = 12'he73;
15'b0000101001111011000 : color = 12'he73;
15'b0000101001111011001 : color = 12'he73;
15'b0000101001111011010 : color = 12'he72;
15'b0000101001111011011 : color = 12'hf10;
15'b0000101001111011100 : color = 12'hf63;
15'b0000101001111011101 : color = 12'he73;
15'b0000101001111011110 : color = 12'he73;
15'b0000101001111011111 : color = 12'he73;
15'b0000101001111100000 : color = 12'he73;
15'b0000101001111100001 : color = 12'he73;
15'b0000101001111100010 : color = 12'he73;
15'b0000101001111100011 : color = 12'hf51;
15'b0000101001111100100 : color = 12'hf10;
15'b0000101001111100101 : color = 12'hf00;
15'b0000101001111100110 : color = 12'hf00;
15'b0000101001111100111 : color = 12'hf00;
15'b0000101001111101000 : color = 12'hf00;
15'b0000101001111101001 : color = 12'hf00;
15'b0000101001111101010 : color = 12'hf00;
15'b0000101001111101011 : color = 12'hf00;
15'b0000101001111101100 : color = 12'hf00;
15'b0000101001111101101 : color = 12'hf00;
15'b0000101001111101110 : color = 12'hf00;
15'b0000101001111101111 : color = 12'hf00;
15'b0000101001111110000 : color = 12'hf00;
15'b0000101001111110001 : color = 12'hf00;
15'b0000101001111110010 : color = 12'hf00;
15'b0000101001111110011 : color = 12'hf42;
15'b0000101001111110100 : color = 12'hf73;
15'b0000101001111110101 : color = 12'he73;
15'b0000101001111110110 : color = 12'he73;
15'b0000101001111110111 : color = 12'he73;
15'b0000101001111111000 : color = 12'he73;
15'b0000101001111111001 : color = 12'he73;
15'b0000101001111111010 : color = 12'he73;
15'b0000101001111111011 : color = 12'he73;
15'b0000101001111111100 : color = 12'he73;
15'b0000101001111111101 : color = 12'he73;
15'b0000101001111111110 : color = 12'he73;
15'b0000101001111111111 : color = 12'he73;
15'b0000101010000000000 : color = 12'he73;
15'b0000101010000000001 : color = 12'he73;
15'b0000101010000000010 : color = 12'he73;
15'b0000101010000000011 : color = 12'he73;
15'b0000101010000000100 : color = 12'he73;
15'b0000101010000000101 : color = 12'he73;
15'b0000101010000000110 : color = 12'he73;
15'b0000101010000000111 : color = 12'he72;
15'b0000101010000001000 : color = 12'hf11;
15'b0000101010000001001 : color = 12'hf73;
15'b0000101010000001010 : color = 12'he73;
15'b0000101010000001011 : color = 12'he73;
15'b0000101010000001100 : color = 12'he73;
15'b0000101010000001101 : color = 12'he73;
15'b0000101010000001110 : color = 12'he73;
15'b0000101010000001111 : color = 12'he73;
15'b0000101010000010000 : color = 12'he73;
15'b0000101010000010001 : color = 12'he73;
15'b0000101010000010010 : color = 12'he62;
15'b0000101010000010011 : color = 12'hf41;
15'b0000101010000010100 : color = 12'hf00;
15'b0000101010000010101 : color = 12'hf10;
15'b0000101010000010110 : color = 12'hf10;
15'b0000101010000010111 : color = 12'hf00;
15'b0000101010000011000 : color = 12'hf00;
15'b0000101010000011001 : color = 12'hf53;
15'b0000101010000011010 : color = 12'he73;
15'b0000101010000011011 : color = 12'he73;
15'b0000101010000011100 : color = 12'he73;
15'b0000101010000011101 : color = 12'he73;
15'b0000101010000011110 : color = 12'he73;
15'b0000101010000011111 : color = 12'he73;
15'b0000101010000100000 : color = 12'he73;
15'b0000101010000100001 : color = 12'he73;
15'b0000101010000100010 : color = 12'he73;
15'b0000101010000100011 : color = 12'he73;
15'b0000101010000100100 : color = 12'he73;
15'b0000101010000100101 : color = 12'he73;
15'b0000101010000100110 : color = 12'he73;
15'b0000101010000100111 : color = 12'he73;
15'b0000101010000101000 : color = 12'he73;
15'b0000101010000101001 : color = 12'he73;
15'b0000101010000101010 : color = 12'he73;
15'b0000101010000101011 : color = 12'he73;
15'b0000101010000101100 : color = 12'he73;
15'b0000101010000101101 : color = 12'he73;
15'b0000101010000101110 : color = 12'he73;
15'b0000101010000101111 : color = 12'he73;
15'b0000101010000110000 : color = 12'he73;
15'b0000101010000110001 : color = 12'he73;
15'b0000101010000110010 : color = 12'he73;
15'b0000101010000110011 : color = 12'he73;
15'b0000101010000110100 : color = 12'he73;
15'b0000101010000110101 : color = 12'he73;
15'b0000101010000110110 : color = 12'he73;
15'b0000101010000110111 : color = 12'he73;
15'b0000101010000111000 : color = 12'hf30;
15'b0000101010000111001 : color = 12'hf00;
15'b0000101010000111010 : color = 12'hf31;
15'b0000101010000111011 : color = 12'hf31;
15'b0000101010000111100 : color = 12'hf31;
15'b0000101010000111101 : color = 12'hf31;
15'b0000101010000111110 : color = 12'hf31;
15'b0000101010000111111 : color = 12'hf31;
15'b0000101010001000000 : color = 12'hf31;
15'b0000101010001000001 : color = 12'hf31;
15'b0000101010001000010 : color = 12'hf31;
15'b0000101010001000011 : color = 12'hf31;
15'b0000101010001000100 : color = 12'hf31;
15'b0000101010001000101 : color = 12'hf00;
15'b0000101010001000110 : color = 12'hf32;
15'b0000101010001000111 : color = 12'he73;
15'b0000101010001001000 : color = 12'he73;
15'b0000101010001001001 : color = 12'he73;
15'b0000101010001001010 : color = 12'he73;
15'b0000101010001001011 : color = 12'he73;
15'b0000101010001001100 : color = 12'he73;
15'b0000101010001001101 : color = 12'he73;
15'b0000101010001001110 : color = 12'he73;
15'b0000101010001001111 : color = 12'he73;
15'b0000101010001010000 : color = 12'he73;
15'b0000101010001010001 : color = 12'he73;
15'b0000101010001010010 : color = 12'he73;
15'b0000101010001010011 : color = 12'he73;
15'b0000101010001010100 : color = 12'he73;
15'b0000101010001010101 : color = 12'he73;
15'b0000101010001010110 : color = 12'he73;
15'b0000101010001010111 : color = 12'he73;
15'b0000101010001011000 : color = 12'he73;
15'b0000101010001011001 : color = 12'he73;
15'b0000101010001011010 : color = 12'he73;
15'b0000101010001011011 : color = 12'he73;
15'b0000101010001011100 : color = 12'he73;
15'b0000101010001011101 : color = 12'he73;
15'b0000101010001011110 : color = 12'he73;
15'b0000101010001011111 : color = 12'he73;
15'b0000101010001100000 : color = 12'he73;
15'b0000101010001100001 : color = 12'he73;
15'b0000101010001100010 : color = 12'he73;
15'b0000101010001100011 : color = 12'he73;
15'b0000101010001100100 : color = 12'he73;
15'b0000101010001100101 : color = 12'he72;
15'b0000101010001100110 : color = 12'hf41;
15'b0000101010001100111 : color = 12'hf31;
15'b0000101010001101000 : color = 12'hf31;
15'b0000101010001101001 : color = 12'hf31;
15'b0000101010001101010 : color = 12'hf31;
15'b0000101010001101011 : color = 12'hf31;
15'b0000101010001101100 : color = 12'hf31;
15'b0000101010001101101 : color = 12'hf31;
15'b0000101010001101110 : color = 12'hf31;
15'b0000101010001101111 : color = 12'hf10;
15'b0000101010001110000 : color = 12'hf10;
15'b0000101010001110001 : color = 12'hf31;
15'b0000101010001110010 : color = 12'hf31;
15'b0000101010001110011 : color = 12'hf31;
15'b0000101010001110100 : color = 12'hf31;
15'b0000101010001110101 : color = 12'hf10;
15'b0000101010001110110 : color = 12'hf00;
15'b0000101010001110111 : color = 12'hf00;
15'b0000101010001111000 : color = 12'hf42;
15'b0000101010001111001 : color = 12'he73;
15'b0000101010001111010 : color = 12'he73;
15'b0000101010001111011 : color = 12'he73;
15'b0000101010001111100 : color = 12'he73;
15'b0000101010001111101 : color = 12'he73;
15'b0000101010001111110 : color = 12'he73;
15'b0000101010001111111 : color = 12'he73;
15'b0000101010010000000 : color = 12'he73;
15'b0000101010010000001 : color = 12'he73;
15'b0000101010010000010 : color = 12'he73;
15'b0000101010010000011 : color = 12'he73;
15'b0000101010010000100 : color = 12'he73;
15'b0000101010010000101 : color = 12'he73;
15'b0000101010010000110 : color = 12'he73;
15'b0000101010010000111 : color = 12'he73;
15'b0000101010010001000 : color = 12'he73;
15'b0000101010010001001 : color = 12'he73;
15'b0000101010010001010 : color = 12'he73;
15'b0000101010010001011 : color = 12'he73;
15'b0000101010010001100 : color = 12'hf40;
15'b0000101010010001101 : color = 12'hf11;
15'b0000101010010001110 : color = 12'hf63;
15'b0000101010010001111 : color = 12'he73;
15'b0000101010010010000 : color = 12'he73;
15'b0000101010010010001 : color = 12'he73;
15'b0000101010010010010 : color = 12'he73;
15'b0000101010010010011 : color = 12'hf51;
15'b0000101010010010100 : color = 12'hf10;
15'b0000101010010010101 : color = 12'hf00;
15'b0000101010010010110 : color = 12'hf10;
15'b0000101010010010111 : color = 12'hf00;
15'b0000101010010011000 : color = 12'hf00;
15'b0000101010010011001 : color = 12'hf53;
15'b0000101010010011010 : color = 12'he73;
15'b0000101010010011011 : color = 12'he73;
15'b0000101010010011100 : color = 12'he73;
15'b0000101010010011101 : color = 12'he73;
15'b0000101010010011110 : color = 12'he73;
15'b0000101010010011111 : color = 12'he73;
15'b0000101010010100000 : color = 12'he72;
15'b0000101010010100001 : color = 12'hf10;
15'b0000101010010100010 : color = 12'hf00;
15'b0000101010010100011 : color = 12'hf63;
15'b0000101010010100100 : color = 12'he73;
15'b0000101010010100101 : color = 12'he73;
15'b0000101010010100110 : color = 12'he73;
15'b0000101010010100111 : color = 12'he73;
15'b0000101010010101000 : color = 12'he73;
15'b0000101010010101001 : color = 12'he73;
15'b0000101010010101010 : color = 12'he73;
15'b0000101010010101011 : color = 12'he73;
15'b0000101010010101100 : color = 12'he73;
15'b0000101010010101101 : color = 12'he73;
15'b0000101010010101110 : color = 12'he73;
15'b0000101010010101111 : color = 12'he73;
15'b0000101010010110000 : color = 12'he73;
15'b0000101010010110001 : color = 12'he73;
15'b0000101010010110010 : color = 12'he73;
15'b0000101010010110011 : color = 12'he73;
15'b0000101010010110100 : color = 12'he73;
15'b0000101010010110101 : color = 12'he73;
15'b0000101010010110110 : color = 12'he73;
15'b0000101010010110111 : color = 12'he73;
15'b0000101010010111000 : color = 12'he73;
15'b0000101010010111001 : color = 12'he73;
15'b0000101010010111010 : color = 12'he73;
15'b0000101010010111011 : color = 12'he73;
15'b0000101010010111100 : color = 12'he73;
15'b0000101010010111101 : color = 12'he73;
15'b0000101010010111110 : color = 12'he73;
15'b0000101010010111111 : color = 12'he73;
15'b0000101010011000000 : color = 12'he72;
15'b0000101010011000001 : color = 12'hf30;
15'b0000101010011000010 : color = 12'hf00;
15'b0000101010011000011 : color = 12'hf63;
15'b0000101010011000100 : color = 12'he73;
15'b0000101010011000101 : color = 12'he73;
15'b0000101010011000110 : color = 12'he73;
15'b0000101010011000111 : color = 12'he73;
15'b0000101010011001000 : color = 12'he73;
15'b0000101010011001001 : color = 12'hf30;
15'b0000101010011001010 : color = 12'hf00;
15'b0000101010011001011 : color = 12'hf42;
15'b0000101010011001100 : color = 12'hf52;
15'b0000101010011001101 : color = 12'hf51;
15'b0000101010011001110 : color = 12'hf10;
15'b0000101010011001111 : color = 12'hf00;
15'b0000101010011010000 : color = 12'hf42;
15'b0000101010011010001 : color = 12'he73;
15'b0000101010011010010 : color = 12'he73;
15'b0000101010011010011 : color = 12'he73;
15'b0000101010011010100 : color = 12'he73;
15'b0000101010011010101 : color = 12'he73;
15'b0000101010011010110 : color = 12'he73;
15'b0000101010011010111 : color = 12'he73;
15'b0000101010011011000 : color = 12'he73;
15'b0000101010011011001 : color = 12'he73;
15'b0000101010011011010 : color = 12'he73;
15'b0000101010011011011 : color = 12'he73;
15'b0000101010011011100 : color = 12'he73;
15'b0000101010011011101 : color = 12'he73;
15'b0000101010011011110 : color = 12'he73;
15'b0000101010011011111 : color = 12'he73;
15'b0000101010011100000 : color = 12'he73;
15'b0000101001100011111 : color = 12'he73;
15'b0000101001100100000 : color = 12'he73;
15'b0000101001100100001 : color = 12'he73;
15'b0000101001100100010 : color = 12'he73;
15'b0000101001100100011 : color = 12'he73;
15'b0000101001100100100 : color = 12'he73;
15'b0000101001100100101 : color = 12'he73;
15'b0000101001100100110 : color = 12'he73;
15'b0000101001100100111 : color = 12'he73;
15'b0000101001100101000 : color = 12'he73;
15'b0000101001100101001 : color = 12'he73;
15'b0000101001100101010 : color = 12'he73;
15'b0000101001100101011 : color = 12'he73;
15'b0000101001100101100 : color = 12'he73;
15'b0000101001100101101 : color = 12'he73;
15'b0000101001100101110 : color = 12'hf51;
15'b0000101001100101111 : color = 12'hf31;
15'b0000101001100110000 : color = 12'hf63;
15'b0000101001100110001 : color = 12'he73;
15'b0000101001100110010 : color = 12'he73;
15'b0000101001100110011 : color = 12'he73;
15'b0000101001100110100 : color = 12'he73;
15'b0000101001100110101 : color = 12'he73;
15'b0000101001100110110 : color = 12'he73;
15'b0000101001100110111 : color = 12'he73;
15'b0000101001100111000 : color = 12'he73;
15'b0000101001100111001 : color = 12'he73;
15'b0000101001100111010 : color = 12'he73;
15'b0000101001100111011 : color = 12'he73;
15'b0000101001100111100 : color = 12'he73;
15'b0000101001100111101 : color = 12'he73;
15'b0000101001100111110 : color = 12'he72;
15'b0000101001100111111 : color = 12'hf63;
15'b0000101001101000000 : color = 12'he73;
15'b0000101001101000001 : color = 12'he73;
15'b0000101001101000010 : color = 12'he73;
15'b0000101001101000011 : color = 12'he73;
15'b0000101001101000100 : color = 12'he73;
15'b0000101001101000101 : color = 12'he73;
15'b0000101001101000110 : color = 12'he73;
15'b0000101001101000111 : color = 12'he73;
15'b0000101001101001000 : color = 12'he73;
15'b0000101001101001001 : color = 12'he73;
15'b0000101001101001010 : color = 12'he73;
15'b0000101001101001011 : color = 12'he73;
15'b0000101001101001100 : color = 12'he73;
15'b0000101001101001101 : color = 12'he73;
15'b0000101001101001110 : color = 12'he73;
15'b0000101001101001111 : color = 12'he73;
15'b0000101001101010000 : color = 12'he73;
15'b0000101001101010001 : color = 12'he73;
15'b0000101001101010010 : color = 12'he73;
15'b0000101001101010011 : color = 12'he73;
15'b0000101001101010100 : color = 12'he73;
15'b0000101001101010101 : color = 12'he73;
15'b0000101001101010110 : color = 12'he73;
15'b0000101001101010111 : color = 12'he73;
15'b0000101001101011000 : color = 12'he73;
15'b0000101001101011001 : color = 12'he73;
15'b0000101001101011010 : color = 12'he73;
15'b0000101001101011011 : color = 12'he73;
15'b0000101001101011100 : color = 12'he73;
15'b0000101001101011101 : color = 12'he73;
15'b0000101001101011110 : color = 12'he73;
15'b0000101001101011111 : color = 12'he73;
15'b0000101001101100000 : color = 12'he73;
15'b0000101001101100001 : color = 12'he73;
15'b0000101001101100010 : color = 12'he73;
15'b0000101001101100011 : color = 12'he73;
15'b0000101001101100100 : color = 12'he73;
15'b0000101001101100101 : color = 12'he73;
15'b0000101001101100110 : color = 12'he73;
15'b0000101001101100111 : color = 12'he73;
15'b0000101001101101000 : color = 12'he73;
15'b0000101001101101001 : color = 12'he73;
15'b0000101001101101010 : color = 12'he73;
15'b0000101001101101011 : color = 12'he73;
15'b0000101001101101100 : color = 12'he73;
15'b0000101001101101101 : color = 12'he73;
15'b0000101001101101110 : color = 12'he73;
15'b0000101001101101111 : color = 12'he73;
15'b0000101001101110000 : color = 12'he73;
15'b0000101001101110001 : color = 12'he73;
15'b0000101001101110010 : color = 12'he73;
15'b0000101001101110011 : color = 12'he73;
15'b0000101001101110100 : color = 12'he73;
15'b0000101001101110101 : color = 12'he73;
15'b0000101001101110110 : color = 12'he73;
15'b0000101001101110111 : color = 12'he73;
15'b0000101001101111000 : color = 12'he73;
15'b0000101001101111001 : color = 12'he73;
15'b0000101001101111010 : color = 12'he73;
15'b0000101001101111011 : color = 12'he73;
15'b0000101001101111100 : color = 12'he73;
15'b0000101001101111101 : color = 12'he73;
15'b0000101001101111110 : color = 12'he73;
15'b0000101001101111111 : color = 12'hf51;
15'b0000101001110000000 : color = 12'hf42;
15'b0000101001110000001 : color = 12'hf73;
15'b0000101001110000010 : color = 12'he73;
15'b0000101001110000011 : color = 12'he73;
15'b0000101001110000100 : color = 12'he73;
15'b0000101001110000101 : color = 12'he73;
15'b0000101001110000110 : color = 12'he73;
15'b0000101001110000111 : color = 12'he73;
15'b0000101001110001000 : color = 12'he73;
15'b0000101001110001001 : color = 12'he73;
15'b0000101001110001010 : color = 12'he73;
15'b0000101001110001011 : color = 12'hf40;
15'b0000101001110001100 : color = 12'hf00;
15'b0000101001110001101 : color = 12'hf53;
15'b0000101001110001110 : color = 12'he73;
15'b0000101001110001111 : color = 12'he73;
15'b0000101001110010000 : color = 12'he73;
15'b0000101001110010001 : color = 12'he73;
15'b0000101001110010010 : color = 12'he73;
15'b0000101001110010011 : color = 12'he73;
15'b0000101001110010100 : color = 12'he73;
15'b0000101001110010101 : color = 12'he73;
15'b0000101001110010110 : color = 12'he73;
15'b0000101001110010111 : color = 12'he73;
15'b0000101001110011000 : color = 12'he73;
15'b0000101001110011001 : color = 12'he73;
15'b0000101001110011010 : color = 12'he73;
15'b0000101001110011011 : color = 12'he73;
15'b0000101001110011100 : color = 12'he73;
15'b0000101001110011101 : color = 12'he73;
15'b0000101001110011110 : color = 12'he73;
15'b0000101001110011111 : color = 12'he73;
15'b0000101001110100000 : color = 12'he73;
15'b0000101001110100001 : color = 12'he73;
15'b0000101001110100010 : color = 12'he73;
15'b0000101001110100011 : color = 12'he73;
15'b0000101001110100100 : color = 12'he73;
15'b0000101001110100101 : color = 12'he73;
15'b0000101001110100110 : color = 12'he73;
15'b0000101001110100111 : color = 12'he73;
15'b0000101001110101000 : color = 12'he73;
15'b0000101001110101001 : color = 12'he73;
15'b0000101001110101010 : color = 12'he73;
15'b0000101001110101011 : color = 12'he73;
15'b0000101001110101100 : color = 12'he61;
15'b0000101001110101101 : color = 12'hf11;
15'b0000101001110101110 : color = 12'hf52;
15'b0000101001110101111 : color = 12'he73;
15'b0000101001110110000 : color = 12'he73;
15'b0000101001110110001 : color = 12'he73;
15'b0000101001110110010 : color = 12'he73;
15'b0000101001110110011 : color = 12'he73;
15'b0000101001110110100 : color = 12'he73;
15'b0000101001110110101 : color = 12'he73;
15'b0000101001110110110 : color = 12'he73;
15'b0000101001110110111 : color = 12'he73;
15'b0000101001110111000 : color = 12'he73;
15'b0000101001110111001 : color = 12'he73;
15'b0000101001110111010 : color = 12'he73;
15'b0000101001110111011 : color = 12'he73;
15'b0000101001110111100 : color = 12'he73;
15'b0000101001110111101 : color = 12'he73;
15'b0000101001110111110 : color = 12'he73;
15'b0000101001110111111 : color = 12'he72;
15'b0000101001111000000 : color = 12'hf40;
15'b0000101001111000001 : color = 12'hf00;
15'b0000101001111000010 : color = 12'hf00;
15'b0000101001111000011 : color = 12'hf32;
15'b0000101001111000100 : color = 12'he73;
15'b0000101001111000101 : color = 12'he73;
15'b0000101001111000110 : color = 12'he73;
15'b0000101001111000111 : color = 12'he73;
15'b0000101001111001000 : color = 12'he73;
15'b0000101001111001001 : color = 12'he73;
15'b0000101001111001010 : color = 12'he73;
15'b0000101001111001011 : color = 12'he73;
15'b0000101001111001100 : color = 12'he73;
15'b0000101001111001101 : color = 12'he73;
15'b0000101001111001110 : color = 12'he73;
15'b0000101001111001111 : color = 12'he73;
15'b0000101001111010000 : color = 12'he73;
15'b0000101001111010001 : color = 12'he73;
15'b0000101001111010010 : color = 12'he73;
15'b0000101001111010011 : color = 12'he73;
15'b0000101001111010100 : color = 12'he73;
15'b0000101001111010101 : color = 12'he73;
15'b0000101001111010110 : color = 12'he73;
15'b0000101001111010111 : color = 12'he73;
15'b0000101001111011000 : color = 12'he73;
15'b0000101001111011001 : color = 12'he73;
15'b0000101001111011010 : color = 12'hf51;
15'b0000101001111011011 : color = 12'hf10;
15'b0000101001111011100 : color = 12'hf11;
15'b0000101001111011101 : color = 12'hf62;
15'b0000101001111011110 : color = 12'he73;
15'b0000101001111011111 : color = 12'he73;
15'b0000101001111100000 : color = 12'he73;
15'b0000101001111100001 : color = 12'he73;
15'b0000101001111100010 : color = 12'he73;
15'b0000101001111100011 : color = 12'he73;
15'b0000101001111100100 : color = 12'he73;
15'b0000101001111100101 : color = 12'he73;
15'b0000101001111100110 : color = 12'he73;
15'b0000101001111100111 : color = 12'he73;
15'b0000101001111101000 : color = 12'he73;
15'b0000101001111101001 : color = 12'he73;
15'b0000101001111101010 : color = 12'hf51;
15'b0000101001111101011 : color = 12'hf10;
15'b0000101001111101100 : color = 12'hf00;
15'b0000101001111101101 : color = 12'hf00;
15'b0000101001111101110 : color = 12'hf00;
15'b0000101001111101111 : color = 12'hf00;
15'b0000101001111110000 : color = 12'hf42;
15'b0000101001111110001 : color = 12'he73;
15'b0000101001111110010 : color = 12'he73;
15'b0000101001111110011 : color = 12'he73;
15'b0000101001111110100 : color = 12'he73;
15'b0000101001111110101 : color = 12'he73;
15'b0000101001111110110 : color = 12'he73;
15'b0000101001111110111 : color = 12'he73;
15'b0000101001111111000 : color = 12'he73;
15'b0000101001111111001 : color = 12'he73;
15'b0000101001111111010 : color = 12'he73;
15'b0000101001111111011 : color = 12'he73;
15'b0000101001111111100 : color = 12'he73;
15'b0000101001111111101 : color = 12'he73;
15'b0000101001111111110 : color = 12'he73;
15'b0000101001111111111 : color = 12'he73;
15'b0000101010000000000 : color = 12'he73;
15'b0000101010000000001 : color = 12'he73;
15'b0000101010000000010 : color = 12'he73;
15'b0000101010000000011 : color = 12'he73;
15'b0000101010000000100 : color = 12'he73;
15'b0000101010000000101 : color = 12'he73;
15'b0000101010000000110 : color = 12'he73;
15'b0000101010000000111 : color = 12'he73;
15'b0000101010000001000 : color = 12'he73;
15'b0000101010000001001 : color = 12'he73;
15'b0000101010000001010 : color = 12'he73;
15'b0000101010000001011 : color = 12'he73;
15'b0000101010000001100 : color = 12'he73;
15'b0000101010000001101 : color = 12'he73;
15'b0000101010000001110 : color = 12'he73;
15'b0000101010000001111 : color = 12'hf62;
15'b0000101010000010000 : color = 12'hf41;
15'b0000101010000010001 : color = 12'hf31;
15'b0000101010000010010 : color = 12'hf10;
15'b0000101010000010011 : color = 12'hf10;
15'b0000101010000010100 : color = 12'hf10;
15'b0000101010000010101 : color = 12'hf00;
15'b0000101010000010110 : color = 12'hf00;
15'b0000101010000010111 : color = 12'hf00;
15'b0000101010000011000 : color = 12'hf00;
15'b0000101010000011001 : color = 12'hf00;
15'b0000101010000011010 : color = 12'hf00;
15'b0000101010000011011 : color = 12'hf11;
15'b0000101010000011100 : color = 12'hf73;
15'b0000101010000011101 : color = 12'he73;
15'b0000101010000011110 : color = 12'he73;
15'b0000101010000011111 : color = 12'he73;
15'b0000101010000100000 : color = 12'he73;
15'b0000101010000100001 : color = 12'he73;
15'b0000101010000100010 : color = 12'he73;
15'b0000101010000100011 : color = 12'he73;
15'b0000101010000100100 : color = 12'he73;
15'b0000101010000100101 : color = 12'he73;
15'b0000101010000100110 : color = 12'he73;
15'b0000101010000100111 : color = 12'he73;
15'b0000101010000101000 : color = 12'he73;
15'b0000101010000101001 : color = 12'he73;
15'b0000101010000101010 : color = 12'he73;
15'b0000101010000101011 : color = 12'he73;
15'b0000101010000101100 : color = 12'he73;
15'b0000101010000101101 : color = 12'he73;
15'b0000101010000101110 : color = 12'he73;
15'b0000101010000101111 : color = 12'he72;
15'b0000101010000110000 : color = 12'hf31;
15'b0000101010000110001 : color = 12'hf63;
15'b0000101010000110010 : color = 12'he73;
15'b0000101010000110011 : color = 12'he73;
15'b0000101010000110100 : color = 12'he73;
15'b0000101010000110101 : color = 12'he73;
15'b0000101010000110110 : color = 12'he73;
15'b0000101010000110111 : color = 12'he73;
15'b0000101010000111000 : color = 12'he73;
15'b0000101010000111001 : color = 12'he73;
15'b0000101010000111010 : color = 12'he73;
15'b0000101010000111011 : color = 12'he73;
15'b0000101010000111100 : color = 12'he73;
15'b0000101010000111101 : color = 12'he72;
15'b0000101010000111110 : color = 12'hf30;
15'b0000101010000111111 : color = 12'hf00;
15'b0000101010001000000 : color = 12'hf00;
15'b0000101010001000001 : color = 12'hf11;
15'b0000101010001000010 : color = 12'hf73;
15'b0000101010001000011 : color = 12'he73;
15'b0000101010001000100 : color = 12'he73;
15'b0000101010001000101 : color = 12'he73;
15'b0000101010001000110 : color = 12'he73;
15'b0000101010001000111 : color = 12'he73;
15'b0000101010001001000 : color = 12'he73;
15'b0000101010001001001 : color = 12'he73;
15'b0000101010001001010 : color = 12'he73;
15'b0000101010001001011 : color = 12'he73;
15'b0000101010001001100 : color = 12'he73;
15'b0000101010001001101 : color = 12'he73;
15'b0000101010001001110 : color = 12'he73;
15'b0000101010001001111 : color = 12'he73;
15'b0000101010001010000 : color = 12'he73;
15'b0000101010001010001 : color = 12'he73;
15'b0000101010001010010 : color = 12'he73;
15'b0000101010001010011 : color = 12'he73;
15'b0000101010001010100 : color = 12'he73;
15'b0000101010001010101 : color = 12'he73;
15'b0000101010001010110 : color = 12'he73;
15'b0000101010001010111 : color = 12'he73;
15'b0000101010001011000 : color = 12'he73;
15'b0000101010001011001 : color = 12'he73;
15'b0000101010001011010 : color = 12'he73;
15'b0000101010001011011 : color = 12'he73;
15'b0000101010001011100 : color = 12'he73;
15'b0000101010001011101 : color = 12'he73;
15'b0000101010001011110 : color = 12'he73;
15'b0000101010001011111 : color = 12'he73;
15'b0000101010001100000 : color = 12'he73;
15'b0000101010001100001 : color = 12'hf30;
15'b0000101010001100010 : color = 12'hf11;
15'b0000101010001100011 : color = 12'hf73;
15'b0000101010001100100 : color = 12'he73;
15'b0000101010001100101 : color = 12'he73;
15'b0000101010001100110 : color = 12'he73;
15'b0000101010001100111 : color = 12'he73;
15'b0000101010001101000 : color = 12'he73;
15'b0000101010001101001 : color = 12'he73;
15'b0000101010001101010 : color = 12'he73;
15'b0000101010001101011 : color = 12'he73;
15'b0000101010001101100 : color = 12'he73;
15'b0000101010001101101 : color = 12'he72;
15'b0000101010001101110 : color = 12'hf10;
15'b0000101010001101111 : color = 12'hf32;
15'b0000101010001110000 : color = 12'he73;
15'b0000101010001110001 : color = 12'he73;
15'b0000101010001110010 : color = 12'he73;
15'b0000101010001110011 : color = 12'he73;
15'b0000101010001110100 : color = 12'he73;
15'b0000101010001110101 : color = 12'he73;
15'b0000101010001110110 : color = 12'he73;
15'b0000101010001110111 : color = 12'he73;
15'b0000101010001111000 : color = 12'he73;
15'b0000101010001111001 : color = 12'he73;
15'b0000101010001111010 : color = 12'he73;
15'b0000101010001111011 : color = 12'he73;
15'b0000101010001111100 : color = 12'he73;
15'b0000101010001111101 : color = 12'he73;
15'b0000101010001111110 : color = 12'he73;
15'b0000101010001111111 : color = 12'he73;
15'b0000101010010000000 : color = 12'he73;
15'b0000101010010000001 : color = 12'he73;
15'b0000101010010000010 : color = 12'he73;
15'b0000101010010000011 : color = 12'he73;
15'b0000101010010000100 : color = 12'he73;
15'b0000101010010000101 : color = 12'he73;
15'b0000101010010000110 : color = 12'he73;
15'b0000101010010000111 : color = 12'he73;
15'b0000101010010001000 : color = 12'he73;
15'b0000101010010001001 : color = 12'he73;
15'b0000101010010001010 : color = 12'he73;
15'b0000101010010001011 : color = 12'he73;
15'b0000101010010001100 : color = 12'he73;
15'b0000101010010001101 : color = 12'he73;
15'b0000101010010001110 : color = 12'he73;
15'b0000101010010001111 : color = 12'he72;
15'b0000101010010010000 : color = 12'hf63;
15'b0000101010010010001 : color = 12'he73;
15'b0000101010010010010 : color = 12'he73;
15'b0000101010010010011 : color = 12'he73;
15'b0000101010010010100 : color = 12'he73;
15'b0000101010010010101 : color = 12'he73;
15'b0000101010010010110 : color = 12'he73;
15'b0000101010010010111 : color = 12'he73;
15'b0000101010010011000 : color = 12'he73;
15'b0000101010010011001 : color = 12'he73;
15'b0000101010010011010 : color = 12'he73;
15'b0000101010010011011 : color = 12'he73;
15'b0000101010010011100 : color = 12'he73;
15'b0000101010010011101 : color = 12'he73;
15'b0000101010010011110 : color = 12'he73;
15'b0000101010010011111 : color = 12'he73;
15'b0000101010010100000 : color = 12'he73;
15'b0000101010010100001 : color = 12'he73;
15'b0000101010010100010 : color = 12'he73;
15'b0000101010010100011 : color = 12'he73;
15'b0000101010010100100 : color = 12'he73;
15'b0000101010010100101 : color = 12'he73;
15'b0000101010010100110 : color = 12'he73;
15'b0000101010010100111 : color = 12'he73;
15'b0000101010010101000 : color = 12'he73;
15'b0000101010010101001 : color = 12'he73;
15'b0000101010010101010 : color = 12'he73;
15'b0000101010010101011 : color = 12'he73;
15'b0000101010010101100 : color = 12'he73;
15'b0000101010010101101 : color = 12'he73;
15'b0000101010010101110 : color = 12'he73;
15'b0000101010010101111 : color = 12'he73;
15'b0000101010010110000 : color = 12'he73;
15'b0000101010010110001 : color = 12'he73;
15'b0000101010010110010 : color = 12'he73;
15'b0000101010010110011 : color = 12'he72;
15'b0000101010010110100 : color = 12'hf31;
15'b0000101010010110101 : color = 12'hf52;
15'b0000101010010110110 : color = 12'he73;
15'b0000101010010110111 : color = 12'he73;
15'b0000101010010111000 : color = 12'he73;
15'b0000101010010111001 : color = 12'he73;
15'b0000101010010111010 : color = 12'he73;
15'b0000101010010111011 : color = 12'he73;
15'b0000101010010111100 : color = 12'he73;
15'b0000101010010111101 : color = 12'he73;
15'b0000101010010111110 : color = 12'he62;
15'b0000101010010111111 : color = 12'hf00;
15'b0000101010011000000 : color = 12'hf00;
15'b0000101010011000001 : color = 12'hf11;
15'b0000101010011000010 : color = 12'hf73;
15'b0000101010011000011 : color = 12'he73;
15'b0000101010011000100 : color = 12'he73;
15'b0000101010011000101 : color = 12'he73;
15'b0000101010011000110 : color = 12'he73;
15'b0000101010011000111 : color = 12'he73;
15'b0000101010011001000 : color = 12'he73;
15'b0000101010011001001 : color = 12'he73;
15'b0000101010011001010 : color = 12'he61;
15'b0000101010011001011 : color = 12'hf32;
15'b0000101010011001100 : color = 12'he73;
15'b0000101010011001101 : color = 12'he73;
15'b0000101010011001110 : color = 12'he73;
15'b0000101010011001111 : color = 12'he73;
15'b0000101010011010000 : color = 12'he73;
15'b0000101010011010001 : color = 12'he73;
15'b0000101010011010010 : color = 12'he73;
15'b0000101010011010011 : color = 12'he73;
15'b0000101010011010100 : color = 12'he73;
15'b0000101010011010101 : color = 12'he73;
15'b0000101010011010110 : color = 12'he73;
15'b0000101010011010111 : color = 12'he73;
15'b0000101010011011000 : color = 12'he73;
15'b0000101010011011001 : color = 12'he73;
15'b0000101010011011010 : color = 12'he73;
15'b0000101010011011011 : color = 12'he73;
15'b0000101010011011100 : color = 12'he73;
15'b0000101010011011101 : color = 12'he73;
15'b0000101010011011110 : color = 12'he73;
15'b0000101010011011111 : color = 12'he73;
15'b0000101010011100000 : color = 12'he73;
15'b0000101010011100001 : color = 12'he73;
15'b0000101010011100010 : color = 12'he73;
15'b0000101010011100011 : color = 12'he73;
15'b0000101010011100100 : color = 12'he73;
15'b0000101010011100101 : color = 12'he73;
15'b0000101010011100110 : color = 12'he73;
15'b0000101010011100111 : color = 12'he73;
15'b0000101010011101000 : color = 12'hf51;
15'b0000101010011101001 : color = 12'hf10;
15'b0000101010011101010 : color = 12'hf32;
15'b0000101010011101011 : color = 12'hf73;
15'b0000101010011101100 : color = 12'he73;
15'b0000101010011101101 : color = 12'he73;
15'b0000101010011101110 : color = 12'he73;
15'b0000101010011101111 : color = 12'he73;
15'b0000101010011110000 : color = 12'he73;
15'b0000101010011110001 : color = 12'he73;
15'b0000101010011110010 : color = 12'he61;
15'b0000101010011110011 : color = 12'hf00;
15'b0000101010011110100 : color = 12'hf00;
15'b0000101010011110101 : color = 12'hf00;
15'b0000101010011110110 : color = 12'hf00;
15'b0000101010011110111 : color = 12'hf00;
15'b0000101010011111000 : color = 12'hf11;
15'b0000101010011111001 : color = 12'hf73;
15'b0000101010011111010 : color = 12'he73;
15'b0000101010011111011 : color = 12'he73;
15'b0000101010011111100 : color = 12'he73;
15'b0000101010011111101 : color = 12'he73;
15'b0000101010011111110 : color = 12'he73;
15'b0000101010011111111 : color = 12'he73;
15'b0000101010100000000 : color = 12'he73;
15'b0000101010100000001 : color = 12'he73;
15'b0000101010100000010 : color = 12'he73;
15'b0000101010100000011 : color = 12'he73;
15'b0000101010100000100 : color = 12'he73;
15'b0000101010100000101 : color = 12'he73;
15'b0000101010100000110 : color = 12'he73;
15'b0000101010100000111 : color = 12'he73;
15'b0000101010100001000 : color = 12'he73;
15'b0000101010100001001 : color = 12'he73;
15'b0000101001101001000 : color = 12'he73;
15'b0000101001101001001 : color = 12'he73;
15'b0000101001101001010 : color = 12'he73;
15'b0000101001101001011 : color = 12'he73;
15'b0000101001101001100 : color = 12'he73;
15'b0000101001101001101 : color = 12'he73;
15'b0000101001101001110 : color = 12'he73;
15'b0000101001101001111 : color = 12'he73;
15'b0000101001101010000 : color = 12'he73;
15'b0000101001101010001 : color = 12'he73;
15'b0000101001101010010 : color = 12'he73;
15'b0000101001101010011 : color = 12'he73;
15'b0000101001101010100 : color = 12'he73;
15'b0000101001101010101 : color = 12'he73;
15'b0000101001101010110 : color = 12'he73;
15'b0000101001101010111 : color = 12'he73;
15'b0000101001101011000 : color = 12'he73;
15'b0000101001101011001 : color = 12'he73;
15'b0000101001101011010 : color = 12'he73;
15'b0000101001101011011 : color = 12'he73;
15'b0000101001101011100 : color = 12'he73;
15'b0000101001101011101 : color = 12'he73;
15'b0000101001101011110 : color = 12'he73;
15'b0000101001101011111 : color = 12'he73;
15'b0000101001101100000 : color = 12'he73;
15'b0000101001101100001 : color = 12'he73;
15'b0000101001101100010 : color = 12'he73;
15'b0000101001101100011 : color = 12'he73;
15'b0000101001101100100 : color = 12'he73;
15'b0000101001101100101 : color = 12'he73;
15'b0000101001101100110 : color = 12'he73;
15'b0000101001101100111 : color = 12'he73;
15'b0000101001101101000 : color = 12'he73;
15'b0000101001101101001 : color = 12'he73;
15'b0000101001101101010 : color = 12'he73;
15'b0000101001101101011 : color = 12'he73;
15'b0000101001101101100 : color = 12'he73;
15'b0000101001101101101 : color = 12'he73;
15'b0000101001101101110 : color = 12'he73;
15'b0000101001101101111 : color = 12'he73;
15'b0000101001101110000 : color = 12'he73;
15'b0000101001101110001 : color = 12'he73;
15'b0000101001101110010 : color = 12'he73;
15'b0000101001101110011 : color = 12'he73;
15'b0000101001101110100 : color = 12'he73;
15'b0000101001101110101 : color = 12'he73;
15'b0000101001101110110 : color = 12'he73;
15'b0000101001101110111 : color = 12'he73;
15'b0000101001101111000 : color = 12'he73;
15'b0000101001101111001 : color = 12'he73;
15'b0000101001101111010 : color = 12'he73;
15'b0000101001101111011 : color = 12'he73;
15'b0000101001101111100 : color = 12'he73;
15'b0000101001101111101 : color = 12'he73;
15'b0000101001101111110 : color = 12'he73;
15'b0000101001101111111 : color = 12'he73;
15'b0000101001110000000 : color = 12'he73;
15'b0000101001110000001 : color = 12'he73;
15'b0000101001110000010 : color = 12'he73;
15'b0000101001110000011 : color = 12'he73;
15'b0000101001110000100 : color = 12'he73;
15'b0000101001110000101 : color = 12'he73;
15'b0000101001110000110 : color = 12'he73;
15'b0000101001110000111 : color = 12'he73;
15'b0000101001110001000 : color = 12'he73;
15'b0000101001110001001 : color = 12'he73;
15'b0000101001110001010 : color = 12'he73;
15'b0000101001110001011 : color = 12'he73;
15'b0000101001110001100 : color = 12'he73;
15'b0000101001110001101 : color = 12'he73;
15'b0000101001110001110 : color = 12'he73;
15'b0000101001110001111 : color = 12'he73;
15'b0000101001110010000 : color = 12'he73;
15'b0000101001110010001 : color = 12'he73;
15'b0000101001110010010 : color = 12'he73;
15'b0000101001110010011 : color = 12'he73;
15'b0000101001110010100 : color = 12'he73;
15'b0000101001110010101 : color = 12'he73;
15'b0000101001110010110 : color = 12'he73;
15'b0000101001110010111 : color = 12'he73;
15'b0000101001110011000 : color = 12'he73;
15'b0000101001110011001 : color = 12'he73;
15'b0000101001110011010 : color = 12'he73;
15'b0000101001110011011 : color = 12'he73;
15'b0000101001110011100 : color = 12'he73;
15'b0000101001110011101 : color = 12'he73;
15'b0000101001110011110 : color = 12'he73;
15'b0000101001110011111 : color = 12'he73;
15'b0000101001110100000 : color = 12'he73;
15'b0000101001110100001 : color = 12'he73;
15'b0000101001110100010 : color = 12'he73;
15'b0000101001110100011 : color = 12'he73;
15'b0000101001110100100 : color = 12'he73;
15'b0000101001110100101 : color = 12'he73;
15'b0000101001110100110 : color = 12'he73;
15'b0000101001110100111 : color = 12'he73;
15'b0000101001110101000 : color = 12'he73;
15'b0000101001110101001 : color = 12'he73;
15'b0000101001110101010 : color = 12'he73;
15'b0000101001110101011 : color = 12'he73;
15'b0000101001110101100 : color = 12'he73;
15'b0000101001110101101 : color = 12'he73;
15'b0000101001110101110 : color = 12'he73;
15'b0000101001110101111 : color = 12'he73;
15'b0000101001110110000 : color = 12'he73;
15'b0000101001110110001 : color = 12'he73;
15'b0000101001110110010 : color = 12'he73;
15'b0000101001110110011 : color = 12'he73;
15'b0000101001110110100 : color = 12'hf41;
15'b0000101001110110101 : color = 12'hf42;
15'b0000101001110110110 : color = 12'hf73;
15'b0000101001110110111 : color = 12'he73;
15'b0000101001110111000 : color = 12'he73;
15'b0000101001110111001 : color = 12'he73;
15'b0000101001110111010 : color = 12'he73;
15'b0000101001110111011 : color = 12'he73;
15'b0000101001110111100 : color = 12'he73;
15'b0000101001110111101 : color = 12'he73;
15'b0000101001110111110 : color = 12'he73;
15'b0000101001110111111 : color = 12'he73;
15'b0000101001111000000 : color = 12'he73;
15'b0000101001111000001 : color = 12'he73;
15'b0000101001111000010 : color = 12'he73;
15'b0000101001111000011 : color = 12'he73;
15'b0000101001111000100 : color = 12'he73;
15'b0000101001111000101 : color = 12'he73;
15'b0000101001111000110 : color = 12'he73;
15'b0000101001111000111 : color = 12'he73;
15'b0000101001111001000 : color = 12'he73;
15'b0000101001111001001 : color = 12'he73;
15'b0000101001111001010 : color = 12'he73;
15'b0000101001111001011 : color = 12'he73;
15'b0000101001111001100 : color = 12'he73;
15'b0000101001111001101 : color = 12'he73;
15'b0000101001111001110 : color = 12'he73;
15'b0000101001111001111 : color = 12'he73;
15'b0000101001111010000 : color = 12'he73;
15'b0000101001111010001 : color = 12'he73;
15'b0000101001111010010 : color = 12'he73;
15'b0000101001111010011 : color = 12'he73;
15'b0000101001111010100 : color = 12'he73;
15'b0000101001111010101 : color = 12'he73;
15'b0000101001111010110 : color = 12'he73;
15'b0000101001111010111 : color = 12'he73;
15'b0000101001111011000 : color = 12'he73;
15'b0000101001111011001 : color = 12'he73;
15'b0000101001111011010 : color = 12'he73;
15'b0000101001111011011 : color = 12'he73;
15'b0000101001111011100 : color = 12'he73;
15'b0000101001111011101 : color = 12'he73;
15'b0000101001111011110 : color = 12'he73;
15'b0000101001111011111 : color = 12'he73;
15'b0000101001111100000 : color = 12'he73;
15'b0000101001111100001 : color = 12'he73;
15'b0000101001111100010 : color = 12'he73;
15'b0000101001111100011 : color = 12'he73;
15'b0000101001111100100 : color = 12'he73;
15'b0000101001111100101 : color = 12'he73;
15'b0000101001111100110 : color = 12'he73;
15'b0000101001111100111 : color = 12'he73;
15'b0000101001111101000 : color = 12'he73;
15'b0000101001111101001 : color = 12'he73;
15'b0000101001111101010 : color = 12'hf30;
15'b0000101001111101011 : color = 12'hf32;
15'b0000101001111101100 : color = 12'hf73;
15'b0000101001111101101 : color = 12'he73;
15'b0000101001111101110 : color = 12'he73;
15'b0000101001111101111 : color = 12'he73;
15'b0000101001111110000 : color = 12'he73;
15'b0000101001111110001 : color = 12'he73;
15'b0000101001111110010 : color = 12'he73;
15'b0000101001111110011 : color = 12'he73;
15'b0000101001111110100 : color = 12'he73;
15'b0000101001111110101 : color = 12'he73;
15'b0000101001111110110 : color = 12'he73;
15'b0000101001111110111 : color = 12'he73;
15'b0000101001111111000 : color = 12'he73;
15'b0000101001111111001 : color = 12'he73;
15'b0000101001111111010 : color = 12'he73;
15'b0000101001111111011 : color = 12'he73;
15'b0000101001111111100 : color = 12'he73;
15'b0000101001111111101 : color = 12'he73;
15'b0000101001111111110 : color = 12'he73;
15'b0000101001111111111 : color = 12'he73;
15'b0000101010000000000 : color = 12'he72;
15'b0000101010000000001 : color = 12'hf31;
15'b0000101010000000010 : color = 12'hf31;
15'b0000101010000000011 : color = 12'hf52;
15'b0000101010000000100 : color = 12'he73;
15'b0000101010000000101 : color = 12'he73;
15'b0000101010000000110 : color = 12'he73;
15'b0000101010000000111 : color = 12'he73;
15'b0000101010000001000 : color = 12'he73;
15'b0000101010000001001 : color = 12'he73;
15'b0000101010000001010 : color = 12'he73;
15'b0000101010000001011 : color = 12'he73;
15'b0000101010000001100 : color = 12'he73;
15'b0000101010000001101 : color = 12'he73;
15'b0000101010000001110 : color = 12'he73;
15'b0000101010000001111 : color = 12'he73;
15'b0000101010000010000 : color = 12'he73;
15'b0000101010000010001 : color = 12'he73;
15'b0000101010000010010 : color = 12'he73;
15'b0000101010000010011 : color = 12'he73;
15'b0000101010000010100 : color = 12'he73;
15'b0000101010000010101 : color = 12'he73;
15'b0000101010000010110 : color = 12'hf62;
15'b0000101010000010111 : color = 12'hf51;
15'b0000101010000011000 : color = 12'hf42;
15'b0000101010000011001 : color = 12'hf73;
15'b0000101010000011010 : color = 12'he73;
15'b0000101010000011011 : color = 12'he73;
15'b0000101010000011100 : color = 12'he73;
15'b0000101010000011101 : color = 12'he73;
15'b0000101010000011110 : color = 12'he73;
15'b0000101010000011111 : color = 12'he73;
15'b0000101010000100000 : color = 12'he73;
15'b0000101010000100001 : color = 12'he73;
15'b0000101010000100010 : color = 12'he73;
15'b0000101010000100011 : color = 12'he73;
15'b0000101010000100100 : color = 12'he73;
15'b0000101010000100101 : color = 12'he73;
15'b0000101010000100110 : color = 12'he73;
15'b0000101010000100111 : color = 12'he73;
15'b0000101010000101000 : color = 12'he73;
15'b0000101010000101001 : color = 12'he73;
15'b0000101010000101010 : color = 12'he73;
15'b0000101010000101011 : color = 12'he73;
15'b0000101010000101100 : color = 12'he73;
15'b0000101010000101101 : color = 12'he73;
15'b0000101010000101110 : color = 12'he73;
15'b0000101010000101111 : color = 12'he73;
15'b0000101010000110000 : color = 12'he73;
15'b0000101010000110001 : color = 12'he73;
15'b0000101010000110010 : color = 12'he73;
15'b0000101010000110011 : color = 12'he73;
15'b0000101010000110100 : color = 12'he73;
15'b0000101010000110101 : color = 12'he73;
15'b0000101010000110110 : color = 12'he73;
15'b0000101010000110111 : color = 12'he73;
15'b0000101010000111000 : color = 12'he73;
15'b0000101010000111001 : color = 12'he73;
15'b0000101010000111010 : color = 12'he73;
15'b0000101010000111011 : color = 12'he73;
15'b0000101010000111100 : color = 12'he73;
15'b0000101010000111101 : color = 12'he73;
15'b0000101010000111110 : color = 12'he73;
15'b0000101010000111111 : color = 12'he73;
15'b0000101010001000000 : color = 12'he73;
15'b0000101010001000001 : color = 12'he73;
15'b0000101010001000010 : color = 12'he73;
15'b0000101010001000011 : color = 12'he73;
15'b0000101010001000100 : color = 12'he73;
15'b0000101010001000101 : color = 12'he73;
15'b0000101010001000110 : color = 12'he73;
15'b0000101010001000111 : color = 12'he73;
15'b0000101010001001000 : color = 12'he73;
15'b0000101010001001001 : color = 12'he73;
15'b0000101010001001010 : color = 12'he73;
15'b0000101010001001011 : color = 12'he73;
15'b0000101010001001100 : color = 12'he73;
15'b0000101010001001101 : color = 12'he73;
15'b0000101010001001110 : color = 12'he73;
15'b0000101010001001111 : color = 12'he73;
15'b0000101010001010000 : color = 12'he73;
15'b0000101010001010001 : color = 12'he73;
15'b0000101010001010010 : color = 12'he73;
15'b0000101010001010011 : color = 12'he73;
15'b0000101010001010100 : color = 12'he73;
15'b0000101010001010101 : color = 12'he73;
15'b0000101010001010110 : color = 12'he73;
15'b0000101010001010111 : color = 12'he73;
15'b0000101010001011000 : color = 12'he72;
15'b0000101010001011001 : color = 12'hf73;
15'b0000101010001011010 : color = 12'he73;
15'b0000101010001011011 : color = 12'he73;
15'b0000101010001011100 : color = 12'he73;
15'b0000101010001011101 : color = 12'he73;
15'b0000101010001011110 : color = 12'he73;
15'b0000101010001011111 : color = 12'he73;
15'b0000101010001100000 : color = 12'he73;
15'b0000101010001100001 : color = 12'he73;
15'b0000101010001100010 : color = 12'he73;
15'b0000101010001100011 : color = 12'he73;
15'b0000101010001100100 : color = 12'he73;
15'b0000101010001100101 : color = 12'he73;
15'b0000101010001100110 : color = 12'he73;
15'b0000101010001100111 : color = 12'he73;
15'b0000101010001101000 : color = 12'hf30;
15'b0000101010001101001 : color = 12'hf31;
15'b0000101010001101010 : color = 12'hf73;
15'b0000101010001101011 : color = 12'he73;
15'b0000101010001101100 : color = 12'he73;
15'b0000101010001101101 : color = 12'he73;
15'b0000101010001101110 : color = 12'he73;
15'b0000101010001101111 : color = 12'he73;
15'b0000101010001110000 : color = 12'he73;
15'b0000101010001110001 : color = 12'he73;
15'b0000101010001110010 : color = 12'he73;
15'b0000101010001110011 : color = 12'he73;
15'b0000101010001110100 : color = 12'he73;
15'b0000101010001110101 : color = 12'he73;
15'b0000101010001110110 : color = 12'he73;
15'b0000101010001110111 : color = 12'he73;
15'b0000101010001111000 : color = 12'he73;
15'b0000101010001111001 : color = 12'he73;
15'b0000101010001111010 : color = 12'he73;
15'b0000101010001111011 : color = 12'he73;
15'b0000101010001111100 : color = 12'he73;
15'b0000101010001111101 : color = 12'he73;
15'b0000101010001111110 : color = 12'he73;
15'b0000101010001111111 : color = 12'he73;
15'b0000101010010000000 : color = 12'he73;
15'b0000101010010000001 : color = 12'he73;
15'b0000101010010000010 : color = 12'he73;
15'b0000101010010000011 : color = 12'he73;
15'b0000101010010000100 : color = 12'he73;
15'b0000101010010000101 : color = 12'he73;
15'b0000101010010000110 : color = 12'he73;
15'b0000101010010000111 : color = 12'he73;
15'b0000101010010001000 : color = 12'he73;
15'b0000101010010001001 : color = 12'he73;
15'b0000101010010001010 : color = 12'hf30;
15'b0000101010010001011 : color = 12'hf32;
15'b0000101010010001100 : color = 12'hf73;
15'b0000101010010001101 : color = 12'he73;
15'b0000101010010001110 : color = 12'he73;
15'b0000101010010001111 : color = 12'he73;
15'b0000101010010010000 : color = 12'he73;
15'b0000101010010010001 : color = 12'he73;
15'b0000101010010010010 : color = 12'he73;
15'b0000101010010010011 : color = 12'he73;
15'b0000101010010010100 : color = 12'he73;
15'b0000101010010010101 : color = 12'he73;
15'b0000101010010010110 : color = 12'he72;
15'b0000101010010010111 : color = 12'hf52;
15'b0000101010010011000 : color = 12'hf73;
15'b0000101010010011001 : color = 12'he73;
15'b0000101010010011010 : color = 12'he73;
15'b0000101010010011011 : color = 12'he73;
15'b0000101010010011100 : color = 12'he73;
15'b0000101010010011101 : color = 12'he73;
15'b0000101010010011110 : color = 12'he73;
15'b0000101010010011111 : color = 12'he73;
15'b0000101010010100000 : color = 12'he73;
15'b0000101010010100001 : color = 12'he73;
15'b0000101010010100010 : color = 12'he73;
15'b0000101010010100011 : color = 12'he73;
15'b0000101010010100100 : color = 12'he73;
15'b0000101010010100101 : color = 12'he73;
15'b0000101010010100110 : color = 12'he73;
15'b0000101010010100111 : color = 12'he73;
15'b0000101010010101000 : color = 12'he73;
15'b0000101010010101001 : color = 12'he73;
15'b0000101010010101010 : color = 12'he73;
15'b0000101010010101011 : color = 12'he73;
15'b0000101010010101100 : color = 12'he73;
15'b0000101010010101101 : color = 12'he73;
15'b0000101010010101110 : color = 12'he73;
15'b0000101010010101111 : color = 12'he73;
15'b0000101010010110000 : color = 12'he73;
15'b0000101010010110001 : color = 12'he73;
15'b0000101010010110010 : color = 12'he73;
15'b0000101010010110011 : color = 12'he73;
15'b0000101010010110100 : color = 12'he73;
15'b0000101010010110101 : color = 12'he73;
15'b0000101010010110110 : color = 12'he73;
15'b0000101010010110111 : color = 12'he73;
15'b0000101010010111000 : color = 12'he73;
15'b0000101010010111001 : color = 12'he73;
15'b0000101010010111010 : color = 12'he73;
15'b0000101010010111011 : color = 12'he73;
15'b0000101010010111100 : color = 12'he73;
15'b0000101010010111101 : color = 12'he73;
15'b0000101010010111110 : color = 12'he73;
15'b0000101010010111111 : color = 12'he73;
15'b0000101010011000000 : color = 12'he73;
15'b0000101010011000001 : color = 12'he73;
15'b0000101010011000010 : color = 12'he73;
15'b0000101010011000011 : color = 12'he73;
15'b0000101010011000100 : color = 12'he73;
15'b0000101010011000101 : color = 12'he73;
15'b0000101010011000110 : color = 12'he73;
15'b0000101010011000111 : color = 12'he73;
15'b0000101010011001000 : color = 12'he73;
15'b0000101010011001001 : color = 12'he73;
15'b0000101010011001010 : color = 12'he73;
15'b0000101010011001011 : color = 12'he73;
15'b0000101010011001100 : color = 12'he73;
15'b0000101010011001101 : color = 12'he73;
15'b0000101010011001110 : color = 12'he73;
15'b0000101010011001111 : color = 12'he73;
15'b0000101010011010000 : color = 12'he73;
15'b0000101010011010001 : color = 12'he73;
15'b0000101010011010010 : color = 12'he73;
15'b0000101010011010011 : color = 12'he73;
15'b0000101010011010100 : color = 12'he73;
15'b0000101010011010101 : color = 12'he73;
15'b0000101010011010110 : color = 12'he73;
15'b0000101010011010111 : color = 12'he73;
15'b0000101010011011000 : color = 12'he73;
15'b0000101010011011001 : color = 12'he73;
15'b0000101010011011010 : color = 12'he73;
15'b0000101010011011011 : color = 12'he73;
15'b0000101010011011100 : color = 12'he73;
15'b0000101010011011101 : color = 12'he73;
15'b0000101010011011110 : color = 12'he73;
15'b0000101010011011111 : color = 12'he73;
15'b0000101010011100000 : color = 12'he73;
15'b0000101010011100001 : color = 12'he73;
15'b0000101010011100010 : color = 12'he73;
15'b0000101010011100011 : color = 12'he73;
15'b0000101010011100100 : color = 12'he73;
15'b0000101010011100101 : color = 12'he73;
15'b0000101010011100110 : color = 12'he73;
15'b0000101010011100111 : color = 12'he73;
15'b0000101010011101000 : color = 12'he51;
15'b0000101010011101001 : color = 12'hf31;
15'b0000101010011101010 : color = 12'hf63;
15'b0000101010011101011 : color = 12'he73;
15'b0000101010011101100 : color = 12'he73;
15'b0000101010011101101 : color = 12'he73;
15'b0000101010011101110 : color = 12'he73;
15'b0000101010011101111 : color = 12'he73;
15'b0000101010011110000 : color = 12'he73;
15'b0000101010011110001 : color = 12'he73;
15'b0000101010011110010 : color = 12'he73;
15'b0000101010011110011 : color = 12'he73;
15'b0000101010011110100 : color = 12'he73;
15'b0000101010011110101 : color = 12'he73;
15'b0000101010011110110 : color = 12'he73;
15'b0000101010011110111 : color = 12'he73;
15'b0000101010011111000 : color = 12'he73;
15'b0000101010011111001 : color = 12'he73;
15'b0000101010011111010 : color = 12'he73;
15'b0000101010011111011 : color = 12'he73;
15'b0000101010011111100 : color = 12'he73;
15'b0000101010011111101 : color = 12'he73;
15'b0000101010011111110 : color = 12'he73;
15'b0000101010011111111 : color = 12'he73;
15'b0000101010100000000 : color = 12'he73;
15'b0000101010100000001 : color = 12'he73;
15'b0000101010100000010 : color = 12'he73;
15'b0000101010100000011 : color = 12'he73;
15'b0000101010100000100 : color = 12'he73;
15'b0000101010100000101 : color = 12'he73;
15'b0000101010100000110 : color = 12'he73;
15'b0000101010100000111 : color = 12'he73;
15'b0000101010100001000 : color = 12'he73;
15'b0000101010100001001 : color = 12'he73;
15'b0000101010100001010 : color = 12'he73;
15'b0000101010100001011 : color = 12'he73;
15'b0000101010100001100 : color = 12'he73;
15'b0000101010100001101 : color = 12'he73;
15'b0000101010100001110 : color = 12'he73;
15'b0000101010100001111 : color = 12'he62;
15'b0000101010100010000 : color = 12'hf31;
15'b0000101010100010001 : color = 12'hf52;
15'b0000101010100010010 : color = 12'hf73;
15'b0000101010100010011 : color = 12'he73;
15'b0000101010100010100 : color = 12'he73;
15'b0000101010100010101 : color = 12'he73;
15'b0000101010100010110 : color = 12'he73;
15'b0000101010100010111 : color = 12'he73;
15'b0000101010100011000 : color = 12'he73;
15'b0000101010100011001 : color = 12'he73;
15'b0000101010100011010 : color = 12'he73;
15'b0000101010100011011 : color = 12'he73;
15'b0000101010100011100 : color = 12'he73;
15'b0000101010100011101 : color = 12'he73;
15'b0000101010100011110 : color = 12'he73;
15'b0000101010100011111 : color = 12'he73;
15'b0000101010100100000 : color = 12'he73;
15'b0000101010100100001 : color = 12'he73;
15'b0000101010100100010 : color = 12'he73;
15'b0000101010100100011 : color = 12'he73;
15'b0000101010100100100 : color = 12'he73;
15'b0000101010100100101 : color = 12'he73;
15'b0000101010100100110 : color = 12'he73;
15'b0000101010100100111 : color = 12'he73;
15'b0000101010100101000 : color = 12'he73;
15'b0000101010100101001 : color = 12'he73;
15'b0000101010100101010 : color = 12'he73;
15'b0000101010100101011 : color = 12'he73;
15'b0000101010100101100 : color = 12'he73;
15'b0000101010100101101 : color = 12'he73;
15'b0000101010100101110 : color = 12'he73;
15'b0000101010100101111 : color = 12'he73;
15'b0000101010100110000 : color = 12'he73;
15'b0000101010100110001 : color = 12'he73;
15'b0000101010100110010 : color = 12'he73;
15'b0000101001101110001 : color = 12'he73;
15'b0000101001101110010 : color = 12'he73;
15'b0000101001101110011 : color = 12'he73;
15'b0000101001101110100 : color = 12'he73;
15'b0000101001101110101 : color = 12'he73;
15'b0000101001101110110 : color = 12'he73;
15'b0000101001101110111 : color = 12'he73;
15'b0000101001101111000 : color = 12'he73;
15'b0000101001101111001 : color = 12'he73;
15'b0000101001101111010 : color = 12'he73;
15'b0000101001101111011 : color = 12'he73;
15'b0000101001101111100 : color = 12'he73;
15'b0000101001101111101 : color = 12'he73;
15'b0000101001101111110 : color = 12'he73;
15'b0000101001101111111 : color = 12'he73;
15'b0000101001110000000 : color = 12'he73;
15'b0000101001110000001 : color = 12'he73;
15'b0000101001110000010 : color = 12'he73;
15'b0000101001110000011 : color = 12'he73;
15'b0000101001110000100 : color = 12'he73;
15'b0000101001110000101 : color = 12'he73;
15'b0000101001110000110 : color = 12'he73;
15'b0000101001110000111 : color = 12'he73;
15'b0000101001110001000 : color = 12'he73;
15'b0000101001110001001 : color = 12'he73;
15'b0000101001110001010 : color = 12'he73;
15'b0000101001110001011 : color = 12'he73;
15'b0000101001110001100 : color = 12'he73;
15'b0000101001110001101 : color = 12'he73;
15'b0000101001110001110 : color = 12'he73;
15'b0000101001110001111 : color = 12'he73;
15'b0000101001110010000 : color = 12'he73;
15'b0000101001110010001 : color = 12'he73;
15'b0000101001110010010 : color = 12'he73;
15'b0000101001110010011 : color = 12'he73;
15'b0000101001110010100 : color = 12'he73;
15'b0000101001110010101 : color = 12'he73;
15'b0000101001110010110 : color = 12'he73;
15'b0000101001110010111 : color = 12'he73;
15'b0000101001110011000 : color = 12'he73;
15'b0000101001110011001 : color = 12'he73;
15'b0000101001110011010 : color = 12'he73;
15'b0000101001110011011 : color = 12'he73;
15'b0000101001110011100 : color = 12'he73;
15'b0000101001110011101 : color = 12'he73;
15'b0000101001110011110 : color = 12'he73;
15'b0000101001110011111 : color = 12'he73;
15'b0000101001110100000 : color = 12'he73;
15'b0000101001110100001 : color = 12'he73;
15'b0000101001110100010 : color = 12'he73;
15'b0000101001110100011 : color = 12'he73;
15'b0000101001110100100 : color = 12'he73;
15'b0000101001110100101 : color = 12'he73;
15'b0000101001110100110 : color = 12'he73;
15'b0000101001110100111 : color = 12'he73;
15'b0000101001110101000 : color = 12'he73;
15'b0000101001110101001 : color = 12'he73;
15'b0000101001110101010 : color = 12'he73;
15'b0000101001110101011 : color = 12'he73;
15'b0000101001110101100 : color = 12'he73;
15'b0000101001110101101 : color = 12'he73;
15'b0000101001110101110 : color = 12'he73;
15'b0000101001110101111 : color = 12'he73;
15'b0000101001110110000 : color = 12'he73;
15'b0000101001110110001 : color = 12'he73;
15'b0000101001110110010 : color = 12'he73;
15'b0000101001110110011 : color = 12'he73;
15'b0000101001110110100 : color = 12'he73;
15'b0000101001110110101 : color = 12'he73;
15'b0000101001110110110 : color = 12'he73;
15'b0000101001110110111 : color = 12'he73;
15'b0000101001110111000 : color = 12'he73;
15'b0000101001110111001 : color = 12'he73;
15'b0000101001110111010 : color = 12'he73;
15'b0000101001110111011 : color = 12'he73;
15'b0000101001110111100 : color = 12'he73;
15'b0000101001110111101 : color = 12'he73;
15'b0000101001110111110 : color = 12'he73;
15'b0000101001110111111 : color = 12'he73;
15'b0000101001111000000 : color = 12'he73;
15'b0000101001111000001 : color = 12'he73;
15'b0000101001111000010 : color = 12'he73;
15'b0000101001111000011 : color = 12'he73;
15'b0000101001111000100 : color = 12'he73;
15'b0000101001111000101 : color = 12'he73;
15'b0000101001111000110 : color = 12'he73;
15'b0000101001111000111 : color = 12'he73;
15'b0000101001111001000 : color = 12'he73;
15'b0000101001111001001 : color = 12'he73;
15'b0000101001111001010 : color = 12'he73;
15'b0000101001111001011 : color = 12'he73;
15'b0000101001111001100 : color = 12'he73;
15'b0000101001111001101 : color = 12'he73;
15'b0000101001111001110 : color = 12'he73;
15'b0000101001111001111 : color = 12'he73;
15'b0000101001111010000 : color = 12'he73;
15'b0000101001111010001 : color = 12'he73;
15'b0000101001111010010 : color = 12'he73;
15'b0000101001111010011 : color = 12'he73;
15'b0000101001111010100 : color = 12'he73;
15'b0000101001111010101 : color = 12'he73;
15'b0000101001111010110 : color = 12'he73;
15'b0000101001111010111 : color = 12'he73;
15'b0000101001111011000 : color = 12'he73;
15'b0000101001111011001 : color = 12'he73;
15'b0000101001111011010 : color = 12'he73;
15'b0000101001111011011 : color = 12'he73;
15'b0000101001111011100 : color = 12'he73;
15'b0000101001111011101 : color = 12'he73;
15'b0000101001111011110 : color = 12'he73;
15'b0000101001111011111 : color = 12'he73;
15'b0000101001111100000 : color = 12'he73;
15'b0000101001111100001 : color = 12'he73;
15'b0000101001111100010 : color = 12'he73;
15'b0000101001111100011 : color = 12'he73;
15'b0000101001111100100 : color = 12'he73;
15'b0000101001111100101 : color = 12'he73;
15'b0000101001111100110 : color = 12'he73;
15'b0000101001111100111 : color = 12'he73;
15'b0000101001111101000 : color = 12'he73;
15'b0000101001111101001 : color = 12'he73;
15'b0000101001111101010 : color = 12'he73;
15'b0000101001111101011 : color = 12'he73;
15'b0000101001111101100 : color = 12'he73;
15'b0000101001111101101 : color = 12'he73;
15'b0000101001111101110 : color = 12'he73;
15'b0000101001111101111 : color = 12'he73;
15'b0000101001111110000 : color = 12'he73;
15'b0000101001111110001 : color = 12'he73;
15'b0000101001111110010 : color = 12'he73;
15'b0000101001111110011 : color = 12'he73;
15'b0000101001111110100 : color = 12'he73;
15'b0000101001111110101 : color = 12'he73;
15'b0000101001111110110 : color = 12'he73;
15'b0000101001111110111 : color = 12'he73;
15'b0000101001111111000 : color = 12'he73;
15'b0000101001111111001 : color = 12'he73;
15'b0000101001111111010 : color = 12'he73;
15'b0000101001111111011 : color = 12'he73;
15'b0000101001111111100 : color = 12'he73;
15'b0000101001111111101 : color = 12'he73;
15'b0000101001111111110 : color = 12'he73;
15'b0000101001111111111 : color = 12'he73;
15'b0000101010000000000 : color = 12'he73;
15'b0000101010000000001 : color = 12'he73;
15'b0000101010000000010 : color = 12'he73;
15'b0000101010000000011 : color = 12'he73;
15'b0000101010000000100 : color = 12'he73;
15'b0000101010000000101 : color = 12'he73;
15'b0000101010000000110 : color = 12'he73;
15'b0000101010000000111 : color = 12'he73;
15'b0000101010000001000 : color = 12'he73;
15'b0000101010000001001 : color = 12'he73;
15'b0000101010000001010 : color = 12'he73;
15'b0000101010000001011 : color = 12'he73;
15'b0000101010000001100 : color = 12'he73;
15'b0000101010000001101 : color = 12'he73;
15'b0000101010000001110 : color = 12'he73;
15'b0000101010000001111 : color = 12'he73;
15'b0000101010000010000 : color = 12'he73;
15'b0000101010000010001 : color = 12'he73;
15'b0000101010000010010 : color = 12'he73;
15'b0000101010000010011 : color = 12'he73;
15'b0000101010000010100 : color = 12'he73;
15'b0000101010000010101 : color = 12'he73;
15'b0000101010000010110 : color = 12'he73;
15'b0000101010000010111 : color = 12'he73;
15'b0000101010000011000 : color = 12'he73;
15'b0000101010000011001 : color = 12'he73;
15'b0000101010000011010 : color = 12'he73;
15'b0000101010000011011 : color = 12'he73;
15'b0000101010000011100 : color = 12'he73;
15'b0000101010000011101 : color = 12'he73;
15'b0000101010000011110 : color = 12'he73;
15'b0000101010000011111 : color = 12'he73;
15'b0000101010000100000 : color = 12'he73;
15'b0000101010000100001 : color = 12'he73;
15'b0000101010000100010 : color = 12'he73;
15'b0000101010000100011 : color = 12'he73;
15'b0000101010000100100 : color = 12'he73;
15'b0000101010000100101 : color = 12'he73;
15'b0000101010000100110 : color = 12'he73;
15'b0000101010000100111 : color = 12'he73;
15'b0000101010000101000 : color = 12'he73;
15'b0000101010000101001 : color = 12'he73;
15'b0000101010000101010 : color = 12'he73;
15'b0000101010000101011 : color = 12'he73;
15'b0000101010000101100 : color = 12'he73;
15'b0000101010000101101 : color = 12'he73;
15'b0000101010000101110 : color = 12'he73;
15'b0000101010000101111 : color = 12'he73;
15'b0000101010000110000 : color = 12'he73;
15'b0000101010000110001 : color = 12'he73;
15'b0000101010000110010 : color = 12'he73;
15'b0000101010000110011 : color = 12'he73;
15'b0000101010000110100 : color = 12'he73;
15'b0000101010000110101 : color = 12'he73;
15'b0000101010000110110 : color = 12'he73;
15'b0000101010000110111 : color = 12'he73;
15'b0000101010000111000 : color = 12'he73;
15'b0000101010000111001 : color = 12'he73;
15'b0000101010000111010 : color = 12'he73;
15'b0000101010000111011 : color = 12'he73;
15'b0000101010000111100 : color = 12'he73;
15'b0000101010000111101 : color = 12'he73;
15'b0000101010000111110 : color = 12'he73;
15'b0000101010000111111 : color = 12'he73;
15'b0000101010001000000 : color = 12'he73;
15'b0000101010001000001 : color = 12'he73;
15'b0000101010001000010 : color = 12'he73;
15'b0000101010001000011 : color = 12'he73;
15'b0000101010001000100 : color = 12'he73;
15'b0000101010001000101 : color = 12'he73;
15'b0000101010001000110 : color = 12'he73;
15'b0000101010001000111 : color = 12'he73;
15'b0000101010001001000 : color = 12'he73;
15'b0000101010001001001 : color = 12'he73;
15'b0000101010001001010 : color = 12'he73;
15'b0000101010001001011 : color = 12'he73;
15'b0000101010001001100 : color = 12'he73;
15'b0000101010001001101 : color = 12'he73;
15'b0000101010001001110 : color = 12'he73;
15'b0000101010001001111 : color = 12'he73;
15'b0000101010001010000 : color = 12'he73;
15'b0000101010001010001 : color = 12'he73;
15'b0000101010001010010 : color = 12'he73;
15'b0000101010001010011 : color = 12'he73;
15'b0000101010001010100 : color = 12'he73;
15'b0000101010001010101 : color = 12'he73;
15'b0000101010001010110 : color = 12'he73;
15'b0000101010001010111 : color = 12'he73;
15'b0000101010001011000 : color = 12'he73;
15'b0000101010001011001 : color = 12'he73;
15'b0000101010001011010 : color = 12'he73;
15'b0000101010001011011 : color = 12'he73;
15'b0000101010001011100 : color = 12'he73;
15'b0000101010001011101 : color = 12'he73;
15'b0000101010001011110 : color = 12'he73;
15'b0000101010001011111 : color = 12'he73;
15'b0000101010001100000 : color = 12'he73;
15'b0000101010001100001 : color = 12'he73;
15'b0000101010001100010 : color = 12'he73;
15'b0000101010001100011 : color = 12'he73;
15'b0000101010001100100 : color = 12'he73;
15'b0000101010001100101 : color = 12'he73;
15'b0000101010001100110 : color = 12'he73;
15'b0000101010001100111 : color = 12'he73;
15'b0000101010001101000 : color = 12'he73;
15'b0000101010001101001 : color = 12'he73;
15'b0000101010001101010 : color = 12'he73;
15'b0000101010001101011 : color = 12'he73;
15'b0000101010001101100 : color = 12'he73;
15'b0000101010001101101 : color = 12'he73;
15'b0000101010001101110 : color = 12'he73;
15'b0000101010001101111 : color = 12'he73;
15'b0000101010001110000 : color = 12'he73;
15'b0000101010001110001 : color = 12'he73;
15'b0000101010001110010 : color = 12'he73;
15'b0000101010001110011 : color = 12'he73;
15'b0000101010001110100 : color = 12'he73;
15'b0000101010001110101 : color = 12'he73;
15'b0000101010001110110 : color = 12'he73;
15'b0000101010001110111 : color = 12'he73;
15'b0000101010001111000 : color = 12'he73;
15'b0000101010001111001 : color = 12'he73;
15'b0000101010001111010 : color = 12'he73;
15'b0000101010001111011 : color = 12'he73;
15'b0000101010001111100 : color = 12'he73;
15'b0000101010001111101 : color = 12'he73;
15'b0000101010001111110 : color = 12'he73;
15'b0000101010001111111 : color = 12'he73;
15'b0000101010010000000 : color = 12'he73;
15'b0000101010010000001 : color = 12'he73;
15'b0000101010010000010 : color = 12'he73;
15'b0000101010010000011 : color = 12'he73;
15'b0000101010010000100 : color = 12'he73;
15'b0000101010010000101 : color = 12'he73;
15'b0000101010010000110 : color = 12'he73;
15'b0000101010010000111 : color = 12'he73;
15'b0000101010010001000 : color = 12'he73;
15'b0000101010010001001 : color = 12'he73;
15'b0000101010010001010 : color = 12'he73;
15'b0000101010010001011 : color = 12'he73;
15'b0000101010010001100 : color = 12'he73;
15'b0000101010010001101 : color = 12'he73;
15'b0000101010010001110 : color = 12'he73;
15'b0000101010010001111 : color = 12'he73;
15'b0000101010010010000 : color = 12'he73;
15'b0000101010010010001 : color = 12'he73;
15'b0000101010010010010 : color = 12'he73;
15'b0000101010010010011 : color = 12'he73;
15'b0000101010010010100 : color = 12'he73;
15'b0000101010010010101 : color = 12'he73;
15'b0000101010010010110 : color = 12'he73;
15'b0000101010010010111 : color = 12'he73;
15'b0000101010010011000 : color = 12'he73;
15'b0000101010010011001 : color = 12'he73;
15'b0000101010010011010 : color = 12'he73;
15'b0000101010010011011 : color = 12'he73;
15'b0000101010010011100 : color = 12'he73;
15'b0000101010010011101 : color = 12'he73;
15'b0000101010010011110 : color = 12'he73;
15'b0000101010010011111 : color = 12'he73;
15'b0000101010010100000 : color = 12'he73;
15'b0000101010010100001 : color = 12'he73;
15'b0000101010010100010 : color = 12'he73;
15'b0000101010010100011 : color = 12'he73;
15'b0000101010010100100 : color = 12'he73;
15'b0000101010010100101 : color = 12'he73;
15'b0000101010010100110 : color = 12'he73;
15'b0000101010010100111 : color = 12'he73;
15'b0000101010010101000 : color = 12'he73;
15'b0000101010010101001 : color = 12'he73;
15'b0000101010010101010 : color = 12'he73;
15'b0000101010010101011 : color = 12'he73;
15'b0000101010010101100 : color = 12'he73;
15'b0000101010010101101 : color = 12'he73;
15'b0000101010010101110 : color = 12'he73;
15'b0000101010010101111 : color = 12'he73;
15'b0000101010010110000 : color = 12'he73;
15'b0000101010010110001 : color = 12'he73;
15'b0000101010010110010 : color = 12'he73;
15'b0000101010010110011 : color = 12'he73;
15'b0000101010010110100 : color = 12'he73;
15'b0000101010010110101 : color = 12'he73;
15'b0000101010010110110 : color = 12'he73;
15'b0000101010010110111 : color = 12'he73;
15'b0000101010010111000 : color = 12'he73;
15'b0000101010010111001 : color = 12'he73;
15'b0000101010010111010 : color = 12'he73;
15'b0000101010010111011 : color = 12'he73;
15'b0000101010010111100 : color = 12'he73;
15'b0000101010010111101 : color = 12'he73;
15'b0000101010010111110 : color = 12'he73;
15'b0000101010010111111 : color = 12'he73;
15'b0000101010011000000 : color = 12'he73;
15'b0000101010011000001 : color = 12'he73;
15'b0000101010011000010 : color = 12'he73;
15'b0000101010011000011 : color = 12'he73;
15'b0000101010011000100 : color = 12'he73;
15'b0000101010011000101 : color = 12'he73;
15'b0000101010011000110 : color = 12'he73;
15'b0000101010011000111 : color = 12'he73;
15'b0000101010011001000 : color = 12'he73;
15'b0000101010011001001 : color = 12'he73;
15'b0000101010011001010 : color = 12'he73;
15'b0000101010011001011 : color = 12'he73;
15'b0000101010011001100 : color = 12'he73;
15'b0000101010011001101 : color = 12'he73;
15'b0000101010011001110 : color = 12'he73;
15'b0000101010011001111 : color = 12'he73;
15'b0000101010011010000 : color = 12'he73;
15'b0000101010011010001 : color = 12'he73;
15'b0000101010011010010 : color = 12'he73;
15'b0000101010011010011 : color = 12'he73;
15'b0000101010011010100 : color = 12'he73;
15'b0000101010011010101 : color = 12'he73;
15'b0000101010011010110 : color = 12'he73;
15'b0000101010011010111 : color = 12'he73;
15'b0000101010011011000 : color = 12'he73;
15'b0000101010011011001 : color = 12'he73;
15'b0000101010011011010 : color = 12'he73;
15'b0000101010011011011 : color = 12'he73;
15'b0000101010011011100 : color = 12'he73;
15'b0000101010011011101 : color = 12'he73;
15'b0000101010011011110 : color = 12'he73;
15'b0000101010011011111 : color = 12'he73;
15'b0000101010011100000 : color = 12'he73;
15'b0000101010011100001 : color = 12'he73;
15'b0000101010011100010 : color = 12'he73;
15'b0000101010011100011 : color = 12'he73;
15'b0000101010011100100 : color = 12'he73;
15'b0000101010011100101 : color = 12'he73;
15'b0000101010011100110 : color = 12'he73;
15'b0000101010011100111 : color = 12'he73;
15'b0000101010011101000 : color = 12'he73;
15'b0000101010011101001 : color = 12'he73;
15'b0000101010011101010 : color = 12'he73;
15'b0000101010011101011 : color = 12'he73;
15'b0000101010011101100 : color = 12'he73;
15'b0000101010011101101 : color = 12'he73;
15'b0000101010011101110 : color = 12'he73;
15'b0000101010011101111 : color = 12'he73;
15'b0000101010011110000 : color = 12'he73;
15'b0000101010011110001 : color = 12'he73;
15'b0000101010011110010 : color = 12'he73;
15'b0000101010011110011 : color = 12'he73;
15'b0000101010011110100 : color = 12'he73;
15'b0000101010011110101 : color = 12'he73;
15'b0000101010011110110 : color = 12'he73;
15'b0000101010011110111 : color = 12'he73;
15'b0000101010011111000 : color = 12'he73;
15'b0000101010011111001 : color = 12'he73;
15'b0000101010011111010 : color = 12'he73;
15'b0000101010011111011 : color = 12'he73;
15'b0000101010011111100 : color = 12'he73;
15'b0000101010011111101 : color = 12'he73;
15'b0000101010011111110 : color = 12'he73;
15'b0000101010011111111 : color = 12'he73;
15'b0000101010100000000 : color = 12'he73;
15'b0000101010100000001 : color = 12'he73;
15'b0000101010100000010 : color = 12'he73;
15'b0000101010100000011 : color = 12'he73;
15'b0000101010100000100 : color = 12'he73;
15'b0000101010100000101 : color = 12'he73;
15'b0000101010100000110 : color = 12'he73;
15'b0000101010100000111 : color = 12'he73;
15'b0000101010100001000 : color = 12'he73;
15'b0000101010100001001 : color = 12'he73;
15'b0000101010100001010 : color = 12'he73;
15'b0000101010100001011 : color = 12'he73;
15'b0000101010100001100 : color = 12'he73;
15'b0000101010100001101 : color = 12'he73;
15'b0000101010100001110 : color = 12'he73;
15'b0000101010100001111 : color = 12'he73;
15'b0000101010100010000 : color = 12'he73;
15'b0000101010100010001 : color = 12'he73;
15'b0000101010100010010 : color = 12'he73;
15'b0000101010100010011 : color = 12'he73;
15'b0000101010100010100 : color = 12'he73;
15'b0000101010100010101 : color = 12'he73;
15'b0000101010100010110 : color = 12'he73;
15'b0000101010100010111 : color = 12'he73;
15'b0000101010100011000 : color = 12'he73;
15'b0000101010100011001 : color = 12'he73;
15'b0000101010100011010 : color = 12'he73;
15'b0000101010100011011 : color = 12'he73;
15'b0000101010100011100 : color = 12'he73;
15'b0000101010100011101 : color = 12'he73;
15'b0000101010100011110 : color = 12'he73;
15'b0000101010100011111 : color = 12'he73;
15'b0000101010100100000 : color = 12'he73;
15'b0000101010100100001 : color = 12'he73;
15'b0000101010100100010 : color = 12'he73;
15'b0000101010100100011 : color = 12'he73;
15'b0000101010100100100 : color = 12'he73;
15'b0000101010100100101 : color = 12'he73;
15'b0000101010100100110 : color = 12'he73;
15'b0000101010100100111 : color = 12'he73;
15'b0000101010100101000 : color = 12'he73;
15'b0000101010100101001 : color = 12'he73;
15'b0000101010100101010 : color = 12'he73;
15'b0000101010100101011 : color = 12'he73;
15'b0000101010100101100 : color = 12'he73;
15'b0000101010100101101 : color = 12'he73;
15'b0000101010100101110 : color = 12'he73;
15'b0000101010100101111 : color = 12'he73;
15'b0000101010100110000 : color = 12'he73;
15'b0000101010100110001 : color = 12'he73;
15'b0000101010100110010 : color = 12'he73;
15'b0000101010100110011 : color = 12'he73;
15'b0000101010100110100 : color = 12'he73;
15'b0000101010100110101 : color = 12'he73;
15'b0000101010100110110 : color = 12'he73;
15'b0000101010100110111 : color = 12'he73;
15'b0000101010100111000 : color = 12'he73;
15'b0000101010100111001 : color = 12'he73;
15'b0000101010100111010 : color = 12'he73;
15'b0000101010100111011 : color = 12'he73;
15'b0000101010100111100 : color = 12'he73;
15'b0000101010100111101 : color = 12'he73;
15'b0000101010100111110 : color = 12'he73;
15'b0000101010100111111 : color = 12'he73;
15'b0000101010101000000 : color = 12'he73;
15'b0000101010101000001 : color = 12'he73;
15'b0000101010101000010 : color = 12'he73;
15'b0000101010101000011 : color = 12'he73;
15'b0000101010101000100 : color = 12'he73;
15'b0000101010101000101 : color = 12'he73;
15'b0000101010101000110 : color = 12'he73;
15'b0000101010101000111 : color = 12'he73;
15'b0000101010101001000 : color = 12'he73;
15'b0000101010101001001 : color = 12'he73;
15'b0000101010101001010 : color = 12'he73;
15'b0000101010101001011 : color = 12'he73;
15'b0000101010101001100 : color = 12'he73;
15'b0000101010101001101 : color = 12'he73;
15'b0000101010101001110 : color = 12'he73;
15'b0000101010101001111 : color = 12'he73;
15'b0000101010101010000 : color = 12'he73;
15'b0000101010101010001 : color = 12'he73;
15'b0000101010101010010 : color = 12'he73;
15'b0000101010101010011 : color = 12'he73;
15'b0000101010101010100 : color = 12'he73;
15'b0000101010101010101 : color = 12'he73;
15'b0000101010101010110 : color = 12'he73;
15'b0000101010101010111 : color = 12'he73;
15'b0000101010101011000 : color = 12'he73;
15'b0000101010101011001 : color = 12'he73;
15'b0000101010101011010 : color = 12'he73;
15'b0000101010101011011 : color = 12'he73;
15'b0000101001110011010 : color = 12'he73;
15'b0000101001110011011 : color = 12'he73;
15'b0000101001110011100 : color = 12'he73;
15'b0000101001110011101 : color = 12'he73;
15'b0000101001110011110 : color = 12'he73;
15'b0000101001110011111 : color = 12'he73;
15'b0000101001110100000 : color = 12'he73;
15'b0000101001110100001 : color = 12'he73;
15'b0000101001110100010 : color = 12'he73;
15'b0000101001110100011 : color = 12'he73;
15'b0000101001110100100 : color = 12'he73;
15'b0000101001110100101 : color = 12'he73;
15'b0000101001110100110 : color = 12'he73;
15'b0000101001110100111 : color = 12'he73;
15'b0000101001110101000 : color = 12'he73;
15'b0000101001110101001 : color = 12'he73;
15'b0000101001110101010 : color = 12'he73;
15'b0000101001110101011 : color = 12'he73;
15'b0000101001110101100 : color = 12'he73;
15'b0000101001110101101 : color = 12'he73;
15'b0000101001110101110 : color = 12'he73;
15'b0000101001110101111 : color = 12'he73;
15'b0000101001110110000 : color = 12'he73;
15'b0000101001110110001 : color = 12'he73;
15'b0000101001110110010 : color = 12'he73;
15'b0000101001110110011 : color = 12'he73;
15'b0000101001110110100 : color = 12'he73;
15'b0000101001110110101 : color = 12'he73;
15'b0000101001110110110 : color = 12'he73;
15'b0000101001110110111 : color = 12'he73;
15'b0000101001110111000 : color = 12'he73;
15'b0000101001110111001 : color = 12'he73;
15'b0000101001110111010 : color = 12'he73;
15'b0000101001110111011 : color = 12'he73;
15'b0000101001110111100 : color = 12'he73;
15'b0000101001110111101 : color = 12'he73;
15'b0000101001110111110 : color = 12'he73;
15'b0000101001110111111 : color = 12'he73;
15'b0000101001111000000 : color = 12'he73;
15'b0000101001111000001 : color = 12'he73;
15'b0000101001111000010 : color = 12'he73;
15'b0000101001111000011 : color = 12'he73;
15'b0000101001111000100 : color = 12'he73;
15'b0000101001111000101 : color = 12'he73;
15'b0000101001111000110 : color = 12'he73;
15'b0000101001111000111 : color = 12'he73;
15'b0000101001111001000 : color = 12'he73;
15'b0000101001111001001 : color = 12'he73;
15'b0000101001111001010 : color = 12'he73;
15'b0000101001111001011 : color = 12'he73;
15'b0000101001111001100 : color = 12'he73;
15'b0000101001111001101 : color = 12'he73;
15'b0000101001111001110 : color = 12'he73;
15'b0000101001111001111 : color = 12'he73;
15'b0000101001111010000 : color = 12'he73;
15'b0000101001111010001 : color = 12'he73;
15'b0000101001111010010 : color = 12'he73;
15'b0000101001111010011 : color = 12'he73;
15'b0000101001111010100 : color = 12'he73;
15'b0000101001111010101 : color = 12'he73;
15'b0000101001111010110 : color = 12'he73;
15'b0000101001111010111 : color = 12'he73;
15'b0000101001111011000 : color = 12'he73;
15'b0000101001111011001 : color = 12'he73;
15'b0000101001111011010 : color = 12'he73;
15'b0000101001111011011 : color = 12'he73;
15'b0000101001111011100 : color = 12'he73;
15'b0000101001111011101 : color = 12'he73;
15'b0000101001111011110 : color = 12'he73;
15'b0000101001111011111 : color = 12'he73;
15'b0000101001111100000 : color = 12'he73;
15'b0000101001111100001 : color = 12'he73;
15'b0000101001111100010 : color = 12'he73;
15'b0000101001111100011 : color = 12'he73;
15'b0000101001111100100 : color = 12'he73;
15'b0000101001111100101 : color = 12'he73;
15'b0000101001111100110 : color = 12'he73;
15'b0000101001111100111 : color = 12'he73;
15'b0000101001111101000 : color = 12'he73;
15'b0000101001111101001 : color = 12'he73;
15'b0000101001111101010 : color = 12'he73;
15'b0000101001111101011 : color = 12'he73;
15'b0000101001111101100 : color = 12'he73;
15'b0000101001111101101 : color = 12'he73;
15'b0000101001111101110 : color = 12'he73;
15'b0000101001111101111 : color = 12'he73;
15'b0000101001111110000 : color = 12'he73;
15'b0000101001111110001 : color = 12'he73;
15'b0000101001111110010 : color = 12'he73;
15'b0000101001111110011 : color = 12'he73;
15'b0000101001111110100 : color = 12'he73;
15'b0000101001111110101 : color = 12'he73;
15'b0000101001111110110 : color = 12'he73;
15'b0000101001111110111 : color = 12'he73;
15'b0000101001111111000 : color = 12'he73;
15'b0000101001111111001 : color = 12'he73;
15'b0000101001111111010 : color = 12'he73;
15'b0000101001111111011 : color = 12'he73;
15'b0000101001111111100 : color = 12'he73;
15'b0000101001111111101 : color = 12'he73;
15'b0000101001111111110 : color = 12'he73;
15'b0000101001111111111 : color = 12'he73;
15'b0000101010000000000 : color = 12'he73;
15'b0000101010000000001 : color = 12'he73;
15'b0000101010000000010 : color = 12'he73;
15'b0000101010000000011 : color = 12'he73;
15'b0000101010000000100 : color = 12'he73;
15'b0000101010000000101 : color = 12'he73;
15'b0000101010000000110 : color = 12'he73;
15'b0000101010000000111 : color = 12'he73;
15'b0000101010000001000 : color = 12'he73;
15'b0000101010000001001 : color = 12'he73;
15'b0000101010000001010 : color = 12'he73;
15'b0000101010000001011 : color = 12'he73;
15'b0000101010000001100 : color = 12'he73;
15'b0000101010000001101 : color = 12'he73;
15'b0000101010000001110 : color = 12'he73;
15'b0000101010000001111 : color = 12'he73;
15'b0000101010000010000 : color = 12'he73;
15'b0000101010000010001 : color = 12'he73;
15'b0000101010000010010 : color = 12'he73;
15'b0000101010000010011 : color = 12'he73;
15'b0000101010000010100 : color = 12'he73;
15'b0000101010000010101 : color = 12'he73;
15'b0000101010000010110 : color = 12'he73;
15'b0000101010000010111 : color = 12'he73;
15'b0000101010000011000 : color = 12'he73;
15'b0000101010000011001 : color = 12'he73;
15'b0000101010000011010 : color = 12'he73;
15'b0000101010000011011 : color = 12'he73;
15'b0000101010000011100 : color = 12'he73;
15'b0000101010000011101 : color = 12'he73;
15'b0000101010000011110 : color = 12'he73;
15'b0000101010000011111 : color = 12'he73;
15'b0000101010000100000 : color = 12'he73;
15'b0000101010000100001 : color = 12'he73;
15'b0000101010000100010 : color = 12'he73;
15'b0000101010000100011 : color = 12'he73;
15'b0000101010000100100 : color = 12'he73;
15'b0000101010000100101 : color = 12'he73;
15'b0000101010000100110 : color = 12'he73;
15'b0000101010000100111 : color = 12'he73;
15'b0000101010000101000 : color = 12'he73;
15'b0000101010000101001 : color = 12'he73;
15'b0000101010000101010 : color = 12'he73;
15'b0000101010000101011 : color = 12'he73;
15'b0000101010000101100 : color = 12'he73;
15'b0000101010000101101 : color = 12'he73;
15'b0000101010000101110 : color = 12'he73;
15'b0000101010000101111 : color = 12'he73;
15'b0000101010000110000 : color = 12'he73;
15'b0000101010000110001 : color = 12'he73;
15'b0000101010000110010 : color = 12'he73;
15'b0000101010000110011 : color = 12'he73;
15'b0000101010000110100 : color = 12'he73;
15'b0000101010000110101 : color = 12'he73;
15'b0000101010000110110 : color = 12'he73;
15'b0000101010000110111 : color = 12'he73;
15'b0000101010000111000 : color = 12'he73;
15'b0000101010000111001 : color = 12'he73;
15'b0000101010000111010 : color = 12'he73;
15'b0000101010000111011 : color = 12'he73;
15'b0000101010000111100 : color = 12'he73;
15'b0000101010000111101 : color = 12'he73;
15'b0000101010000111110 : color = 12'he73;
15'b0000101010000111111 : color = 12'he73;
15'b0000101010001000000 : color = 12'he73;
15'b0000101010001000001 : color = 12'he73;
15'b0000101010001000010 : color = 12'he73;
15'b0000101010001000011 : color = 12'he73;
15'b0000101010001000100 : color = 12'he73;
15'b0000101010001000101 : color = 12'he73;
15'b0000101010001000110 : color = 12'he73;
15'b0000101010001000111 : color = 12'he73;
15'b0000101010001001000 : color = 12'he73;
15'b0000101010001001001 : color = 12'he73;
15'b0000101010001001010 : color = 12'he73;
15'b0000101010001001011 : color = 12'he73;
15'b0000101010001001100 : color = 12'he73;
15'b0000101010001001101 : color = 12'he73;
15'b0000101010001001110 : color = 12'he73;
15'b0000101010001001111 : color = 12'he73;
15'b0000101010001010000 : color = 12'he73;
15'b0000101010001010001 : color = 12'he73;
15'b0000101010001010010 : color = 12'he73;
15'b0000101010001010011 : color = 12'he73;
15'b0000101010001010100 : color = 12'he73;
15'b0000101010001010101 : color = 12'he73;
15'b0000101010001010110 : color = 12'he73;
15'b0000101010001010111 : color = 12'he73;
15'b0000101010001011000 : color = 12'he73;
15'b0000101010001011001 : color = 12'he73;
15'b0000101010001011010 : color = 12'he73;
15'b0000101010001011011 : color = 12'he73;
15'b0000101010001011100 : color = 12'he73;
15'b0000101010001011101 : color = 12'he73;
15'b0000101010001011110 : color = 12'he73;
15'b0000101010001011111 : color = 12'he73;
15'b0000101010001100000 : color = 12'he73;
15'b0000101010001100001 : color = 12'he73;
15'b0000101010001100010 : color = 12'he73;
15'b0000101010001100011 : color = 12'he73;
15'b0000101010001100100 : color = 12'he73;
15'b0000101010001100101 : color = 12'he73;
15'b0000101010001100110 : color = 12'he73;
15'b0000101010001100111 : color = 12'he73;
15'b0000101010001101000 : color = 12'he73;
15'b0000101010001101001 : color = 12'he73;
15'b0000101010001101010 : color = 12'he73;
15'b0000101010001101011 : color = 12'he73;
15'b0000101010001101100 : color = 12'he73;
15'b0000101010001101101 : color = 12'he73;
15'b0000101010001101110 : color = 12'he73;
15'b0000101010001101111 : color = 12'he73;
15'b0000101010001110000 : color = 12'he73;
15'b0000101010001110001 : color = 12'he73;
15'b0000101010001110010 : color = 12'he73;
15'b0000101010001110011 : color = 12'he73;
15'b0000101010001110100 : color = 12'he73;
15'b0000101010001110101 : color = 12'he73;
15'b0000101010001110110 : color = 12'he73;
15'b0000101010001110111 : color = 12'he73;
15'b0000101010001111000 : color = 12'he73;
15'b0000101010001111001 : color = 12'he73;
15'b0000101010001111010 : color = 12'he73;
15'b0000101010001111011 : color = 12'he73;
15'b0000101010001111100 : color = 12'he73;
15'b0000101010001111101 : color = 12'he73;
15'b0000101010001111110 : color = 12'he73;
15'b0000101010001111111 : color = 12'he73;
15'b0000101010010000000 : color = 12'he73;
15'b0000101010010000001 : color = 12'he73;
15'b0000101010010000010 : color = 12'he73;
15'b0000101010010000011 : color = 12'he73;
15'b0000101010010000100 : color = 12'he73;
15'b0000101010010000101 : color = 12'he73;
15'b0000101010010000110 : color = 12'he73;
15'b0000101010010000111 : color = 12'he73;
15'b0000101010010001000 : color = 12'he73;
15'b0000101010010001001 : color = 12'he73;
15'b0000101010010001010 : color = 12'he73;
15'b0000101010010001011 : color = 12'he73;
15'b0000101010010001100 : color = 12'he73;
15'b0000101010010001101 : color = 12'he73;
15'b0000101010010001110 : color = 12'he73;
15'b0000101010010001111 : color = 12'he73;
15'b0000101010010010000 : color = 12'he73;
15'b0000101010010010001 : color = 12'he73;
15'b0000101010010010010 : color = 12'he73;
15'b0000101010010010011 : color = 12'he73;
15'b0000101010010010100 : color = 12'he73;
15'b0000101010010010101 : color = 12'he73;
15'b0000101010010010110 : color = 12'he73;
15'b0000101010010010111 : color = 12'he73;
15'b0000101010010011000 : color = 12'he73;
15'b0000101010010011001 : color = 12'he73;
15'b0000101010010011010 : color = 12'he73;
15'b0000101010010011011 : color = 12'he73;
15'b0000101010010011100 : color = 12'he73;
15'b0000101010010011101 : color = 12'he73;
15'b0000101010010011110 : color = 12'he73;
15'b0000101010010011111 : color = 12'he73;
15'b0000101010010100000 : color = 12'he73;
15'b0000101010010100001 : color = 12'he73;
15'b0000101010010100010 : color = 12'he73;
15'b0000101010010100011 : color = 12'he73;
15'b0000101010010100100 : color = 12'he73;
15'b0000101010010100101 : color = 12'he73;
15'b0000101010010100110 : color = 12'he73;
15'b0000101010010100111 : color = 12'he73;
15'b0000101010010101000 : color = 12'he73;
15'b0000101010010101001 : color = 12'he73;
15'b0000101010010101010 : color = 12'he73;
15'b0000101010010101011 : color = 12'he73;
15'b0000101010010101100 : color = 12'he73;
15'b0000101010010101101 : color = 12'he73;
15'b0000101010010101110 : color = 12'he73;
15'b0000101010010101111 : color = 12'he73;
15'b0000101010010110000 : color = 12'he73;
15'b0000101010010110001 : color = 12'he73;
15'b0000101010010110010 : color = 12'he73;
15'b0000101010010110011 : color = 12'he73;
15'b0000101010010110100 : color = 12'he73;
15'b0000101010010110101 : color = 12'he73;
15'b0000101010010110110 : color = 12'he73;
15'b0000101010010110111 : color = 12'he73;
15'b0000101010010111000 : color = 12'he73;
15'b0000101010010111001 : color = 12'he73;
15'b0000101010010111010 : color = 12'he73;
15'b0000101010010111011 : color = 12'he73;
15'b0000101010010111100 : color = 12'he73;
15'b0000101010010111101 : color = 12'he73;
15'b0000101010010111110 : color = 12'he73;
15'b0000101010010111111 : color = 12'he73;
15'b0000101010011000000 : color = 12'he73;
15'b0000101010011000001 : color = 12'he73;
15'b0000101010011000010 : color = 12'he73;
15'b0000101010011000011 : color = 12'he73;
15'b0000101010011000100 : color = 12'he73;
15'b0000101010011000101 : color = 12'he73;
15'b0000101010011000110 : color = 12'he73;
15'b0000101010011000111 : color = 12'he73;
15'b0000101010011001000 : color = 12'he73;
15'b0000101010011001001 : color = 12'he73;
15'b0000101010011001010 : color = 12'he73;
15'b0000101010011001011 : color = 12'he73;
15'b0000101010011001100 : color = 12'he73;
15'b0000101010011001101 : color = 12'he73;
15'b0000101010011001110 : color = 12'he73;
15'b0000101010011001111 : color = 12'he73;
15'b0000101010011010000 : color = 12'he73;
15'b0000101010011010001 : color = 12'he73;
15'b0000101010011010010 : color = 12'he73;
15'b0000101010011010011 : color = 12'he73;
15'b0000101010011010100 : color = 12'he73;
15'b0000101010011010101 : color = 12'he73;
15'b0000101010011010110 : color = 12'he73;
15'b0000101010011010111 : color = 12'he73;
15'b0000101010011011000 : color = 12'he73;
15'b0000101010011011001 : color = 12'he73;
15'b0000101010011011010 : color = 12'he73;
15'b0000101010011011011 : color = 12'he73;
15'b0000101010011011100 : color = 12'he73;
15'b0000101010011011101 : color = 12'he73;
15'b0000101010011011110 : color = 12'he73;
15'b0000101010011011111 : color = 12'he73;
15'b0000101010011100000 : color = 12'he73;
15'b0000101010011100001 : color = 12'he73;
15'b0000101010011100010 : color = 12'he73;
15'b0000101010011100011 : color = 12'he73;
15'b0000101010011100100 : color = 12'he73;
15'b0000101010011100101 : color = 12'he73;
15'b0000101010011100110 : color = 12'he73;
15'b0000101010011100111 : color = 12'he73;
15'b0000101010011101000 : color = 12'he73;
15'b0000101010011101001 : color = 12'he73;
15'b0000101010011101010 : color = 12'he73;
15'b0000101010011101011 : color = 12'he73;
15'b0000101010011101100 : color = 12'he73;
15'b0000101010011101101 : color = 12'he73;
15'b0000101010011101110 : color = 12'he73;
15'b0000101010011101111 : color = 12'he73;
15'b0000101010011110000 : color = 12'he73;
15'b0000101010011110001 : color = 12'he73;
15'b0000101010011110010 : color = 12'he73;
15'b0000101010011110011 : color = 12'he73;
15'b0000101010011110100 : color = 12'he73;
15'b0000101010011110101 : color = 12'he73;
15'b0000101010011110110 : color = 12'he73;
15'b0000101010011110111 : color = 12'he73;
15'b0000101010011111000 : color = 12'he73;
15'b0000101010011111001 : color = 12'he73;
15'b0000101010011111010 : color = 12'he73;
15'b0000101010011111011 : color = 12'he73;
15'b0000101010011111100 : color = 12'he73;
15'b0000101010011111101 : color = 12'he73;
15'b0000101010011111110 : color = 12'he73;
15'b0000101010011111111 : color = 12'he73;
15'b0000101010100000000 : color = 12'he73;
15'b0000101010100000001 : color = 12'he73;
15'b0000101010100000010 : color = 12'he73;
15'b0000101010100000011 : color = 12'he73;
15'b0000101010100000100 : color = 12'he73;
15'b0000101010100000101 : color = 12'he73;
15'b0000101010100000110 : color = 12'he73;
15'b0000101010100000111 : color = 12'he73;
15'b0000101010100001000 : color = 12'he73;
15'b0000101010100001001 : color = 12'he73;
15'b0000101010100001010 : color = 12'he73;
15'b0000101010100001011 : color = 12'he73;
15'b0000101010100001100 : color = 12'he73;
15'b0000101010100001101 : color = 12'he73;
15'b0000101010100001110 : color = 12'he73;
15'b0000101010100001111 : color = 12'he73;
15'b0000101010100010000 : color = 12'he73;
15'b0000101010100010001 : color = 12'he73;
15'b0000101010100010010 : color = 12'he73;
15'b0000101010100010011 : color = 12'he73;
15'b0000101010100010100 : color = 12'he73;
15'b0000101010100010101 : color = 12'he73;
15'b0000101010100010110 : color = 12'he73;
15'b0000101010100010111 : color = 12'he73;
15'b0000101010100011000 : color = 12'he73;
15'b0000101010100011001 : color = 12'he73;
15'b0000101010100011010 : color = 12'he73;
15'b0000101010100011011 : color = 12'he73;
15'b0000101010100011100 : color = 12'he73;
15'b0000101010100011101 : color = 12'he73;
15'b0000101010100011110 : color = 12'he73;
15'b0000101010100011111 : color = 12'he73;
15'b0000101010100100000 : color = 12'he73;
15'b0000101010100100001 : color = 12'he73;
15'b0000101010100100010 : color = 12'he73;
15'b0000101010100100011 : color = 12'he73;
15'b0000101010100100100 : color = 12'he73;
15'b0000101010100100101 : color = 12'he73;
15'b0000101010100100110 : color = 12'he73;
15'b0000101010100100111 : color = 12'he73;
15'b0000101010100101000 : color = 12'he73;
15'b0000101010100101001 : color = 12'he73;
15'b0000101010100101010 : color = 12'he73;
15'b0000101010100101011 : color = 12'he73;
15'b0000101010100101100 : color = 12'he73;
15'b0000101010100101101 : color = 12'he73;
15'b0000101010100101110 : color = 12'he73;
15'b0000101010100101111 : color = 12'he73;
15'b0000101010100110000 : color = 12'he73;
15'b0000101010100110001 : color = 12'he73;
15'b0000101010100110010 : color = 12'he73;
15'b0000101010100110011 : color = 12'he73;
15'b0000101010100110100 : color = 12'he73;
15'b0000101010100110101 : color = 12'he73;
15'b0000101010100110110 : color = 12'he73;
15'b0000101010100110111 : color = 12'he73;
15'b0000101010100111000 : color = 12'he73;
15'b0000101010100111001 : color = 12'he73;
15'b0000101010100111010 : color = 12'he73;
15'b0000101010100111011 : color = 12'he73;
15'b0000101010100111100 : color = 12'he73;
15'b0000101010100111101 : color = 12'he73;
15'b0000101010100111110 : color = 12'he73;
15'b0000101010100111111 : color = 12'he73;
15'b0000101010101000000 : color = 12'he73;
15'b0000101010101000001 : color = 12'he73;
15'b0000101010101000010 : color = 12'he73;
15'b0000101010101000011 : color = 12'he73;
15'b0000101010101000100 : color = 12'he73;
15'b0000101010101000101 : color = 12'he73;
15'b0000101010101000110 : color = 12'he73;
15'b0000101010101000111 : color = 12'he73;
15'b0000101010101001000 : color = 12'he73;
15'b0000101010101001001 : color = 12'he73;
15'b0000101010101001010 : color = 12'he73;
15'b0000101010101001011 : color = 12'he73;
15'b0000101010101001100 : color = 12'he73;
15'b0000101010101001101 : color = 12'he73;
15'b0000101010101001110 : color = 12'he73;
15'b0000101010101001111 : color = 12'he73;
15'b0000101010101010000 : color = 12'he73;
15'b0000101010101010001 : color = 12'he73;
15'b0000101010101010010 : color = 12'he73;
15'b0000101010101010011 : color = 12'he73;
15'b0000101010101010100 : color = 12'he73;
15'b0000101010101010101 : color = 12'he73;
15'b0000101010101010110 : color = 12'he73;
15'b0000101010101010111 : color = 12'he73;
15'b0000101010101011000 : color = 12'he73;
15'b0000101010101011001 : color = 12'he73;
15'b0000101010101011010 : color = 12'he73;
15'b0000101010101011011 : color = 12'he73;
15'b0000101010101011100 : color = 12'he73;
15'b0000101010101011101 : color = 12'he73;
15'b0000101010101011110 : color = 12'he73;
15'b0000101010101011111 : color = 12'he73;
15'b0000101010101100000 : color = 12'he73;
15'b0000101010101100001 : color = 12'he73;
15'b0000101010101100010 : color = 12'he73;
15'b0000101010101100011 : color = 12'he73;
15'b0000101010101100100 : color = 12'he73;
15'b0000101010101100101 : color = 12'he73;
15'b0000101010101100110 : color = 12'he73;
15'b0000101010101100111 : color = 12'he73;
15'b0000101010101101000 : color = 12'he73;
15'b0000101010101101001 : color = 12'he73;
15'b0000101010101101010 : color = 12'he73;
15'b0000101010101101011 : color = 12'he73;
15'b0000101010101101100 : color = 12'he73;
15'b0000101010101101101 : color = 12'he73;
15'b0000101010101101110 : color = 12'he73;
15'b0000101010101101111 : color = 12'he73;
15'b0000101010101110000 : color = 12'he73;
15'b0000101010101110001 : color = 12'he73;
15'b0000101010101110010 : color = 12'he73;
15'b0000101010101110011 : color = 12'he73;
15'b0000101010101110100 : color = 12'he73;
15'b0000101010101110101 : color = 12'he73;
15'b0000101010101110110 : color = 12'he73;
15'b0000101010101110111 : color = 12'he73;
15'b0000101010101111000 : color = 12'he73;
15'b0000101010101111001 : color = 12'he73;
15'b0000101010101111010 : color = 12'he73;
15'b0000101010101111011 : color = 12'he73;
15'b0000101010101111100 : color = 12'he73;
15'b0000101010101111101 : color = 12'he73;
15'b0000101010101111110 : color = 12'he73;
15'b0000101010101111111 : color = 12'he73;
15'b0000101010110000000 : color = 12'he73;
15'b0000101010110000001 : color = 12'he73;
15'b0000101010110000010 : color = 12'he73;
15'b0000101010110000011 : color = 12'he73;
15'b0000101010110000100 : color = 12'he73;
15'b0000101001111000011 : color = 12'he73;
15'b0000101001111000100 : color = 12'he73;
15'b0000101001111000101 : color = 12'he73;
15'b0000101001111000110 : color = 12'he73;
15'b0000101001111000111 : color = 12'he73;
15'b0000101001111001000 : color = 12'he73;
15'b0000101001111001001 : color = 12'he73;
15'b0000101001111001010 : color = 12'he73;
15'b0000101001111001011 : color = 12'he73;
15'b0000101001111001100 : color = 12'he73;
15'b0000101001111001101 : color = 12'he73;
15'b0000101001111001110 : color = 12'he73;
15'b0000101001111001111 : color = 12'he73;
15'b0000101001111010000 : color = 12'he73;
15'b0000101001111010001 : color = 12'he73;
15'b0000101001111010010 : color = 12'he73;
15'b0000101001111010011 : color = 12'he73;
15'b0000101001111010100 : color = 12'he73;
15'b0000101001111010101 : color = 12'he73;
15'b0000101001111010110 : color = 12'he73;
15'b0000101001111010111 : color = 12'he73;
15'b0000101001111011000 : color = 12'he73;
15'b0000101001111011001 : color = 12'he73;
15'b0000101001111011010 : color = 12'he73;
15'b0000101001111011011 : color = 12'he73;
15'b0000101001111011100 : color = 12'he73;
15'b0000101001111011101 : color = 12'he73;
15'b0000101001111011110 : color = 12'he73;
15'b0000101001111011111 : color = 12'he73;
15'b0000101001111100000 : color = 12'he73;
15'b0000101001111100001 : color = 12'he73;
15'b0000101001111100010 : color = 12'he73;
15'b0000101001111100011 : color = 12'he73;
15'b0000101001111100100 : color = 12'he73;
15'b0000101001111100101 : color = 12'he73;
15'b0000101001111100110 : color = 12'he73;
15'b0000101001111100111 : color = 12'he73;
15'b0000101001111101000 : color = 12'he73;
15'b0000101001111101001 : color = 12'he73;
15'b0000101001111101010 : color = 12'he73;
15'b0000101001111101011 : color = 12'he73;
15'b0000101001111101100 : color = 12'he73;
15'b0000101001111101101 : color = 12'he73;
15'b0000101001111101110 : color = 12'he73;
15'b0000101001111101111 : color = 12'he73;
15'b0000101001111110000 : color = 12'he73;
15'b0000101001111110001 : color = 12'he73;
15'b0000101001111110010 : color = 12'he73;
15'b0000101001111110011 : color = 12'he73;
15'b0000101001111110100 : color = 12'he73;
15'b0000101001111110101 : color = 12'he73;
15'b0000101001111110110 : color = 12'he73;
15'b0000101001111110111 : color = 12'he73;
15'b0000101001111111000 : color = 12'he73;
15'b0000101001111111001 : color = 12'he73;
15'b0000101001111111010 : color = 12'he73;
15'b0000101001111111011 : color = 12'he73;
15'b0000101001111111100 : color = 12'he73;
15'b0000101001111111101 : color = 12'he73;
15'b0000101001111111110 : color = 12'he73;
15'b0000101001111111111 : color = 12'he73;
15'b0000101010000000000 : color = 12'he73;
15'b0000101010000000001 : color = 12'he73;
15'b0000101010000000010 : color = 12'he73;
15'b0000101010000000011 : color = 12'he73;
15'b0000101010000000100 : color = 12'he73;
15'b0000101010000000101 : color = 12'he73;
15'b0000101010000000110 : color = 12'he73;
15'b0000101010000000111 : color = 12'he73;
15'b0000101010000001000 : color = 12'he73;
15'b0000101010000001001 : color = 12'he73;
15'b0000101010000001010 : color = 12'he73;
15'b0000101010000001011 : color = 12'he73;
15'b0000101010000001100 : color = 12'he73;
15'b0000101010000001101 : color = 12'he73;
15'b0000101010000001110 : color = 12'he73;
15'b0000101010000001111 : color = 12'he73;
15'b0000101010000010000 : color = 12'he73;
15'b0000101010000010001 : color = 12'he73;
15'b0000101010000010010 : color = 12'he73;
15'b0000101010000010011 : color = 12'he73;
15'b0000101010000010100 : color = 12'he73;
15'b0000101010000010101 : color = 12'he73;
15'b0000101010000010110 : color = 12'he73;
15'b0000101010000010111 : color = 12'he73;
15'b0000101010000011000 : color = 12'he73;
15'b0000101010000011001 : color = 12'he73;
15'b0000101010000011010 : color = 12'he73;
15'b0000101010000011011 : color = 12'he73;
15'b0000101010000011100 : color = 12'he73;
15'b0000101010000011101 : color = 12'he73;
15'b0000101010000011110 : color = 12'he73;
15'b0000101010000011111 : color = 12'he73;
15'b0000101010000100000 : color = 12'he73;
15'b0000101010000100001 : color = 12'he73;
15'b0000101010000100010 : color = 12'he73;
15'b0000101010000100011 : color = 12'he73;
15'b0000101010000100100 : color = 12'he73;
15'b0000101010000100101 : color = 12'he73;
15'b0000101010000100110 : color = 12'he73;
15'b0000101010000100111 : color = 12'he73;
15'b0000101010000101000 : color = 12'he73;
15'b0000101010000101001 : color = 12'he73;
15'b0000101010000101010 : color = 12'he73;
15'b0000101010000101011 : color = 12'he73;
15'b0000101010000101100 : color = 12'he73;
15'b0000101010000101101 : color = 12'he73;
15'b0000101010000101110 : color = 12'he73;
15'b0000101010000101111 : color = 12'he73;
15'b0000101010000110000 : color = 12'he73;
15'b0000101010000110001 : color = 12'he73;
15'b0000101010000110010 : color = 12'he73;
15'b0000101010000110011 : color = 12'he73;
15'b0000101010000110100 : color = 12'he73;
15'b0000101010000110101 : color = 12'he73;
15'b0000101010000110110 : color = 12'he73;
15'b0000101010000110111 : color = 12'he73;
15'b0000101010000111000 : color = 12'he73;
15'b0000101010000111001 : color = 12'he73;
15'b0000101010000111010 : color = 12'he73;
15'b0000101010000111011 : color = 12'he73;
15'b0000101010000111100 : color = 12'he73;
15'b0000101010000111101 : color = 12'he73;
15'b0000101010000111110 : color = 12'he73;
15'b0000101010000111111 : color = 12'he73;
15'b0000101010001000000 : color = 12'he73;
15'b0000101010001000001 : color = 12'he73;
15'b0000101010001000010 : color = 12'he73;
15'b0000101010001000011 : color = 12'he73;
15'b0000101010001000100 : color = 12'he73;
15'b0000101010001000101 : color = 12'he73;
15'b0000101010001000110 : color = 12'he73;
15'b0000101010001000111 : color = 12'he73;
15'b0000101010001001000 : color = 12'he73;
15'b0000101010001001001 : color = 12'he73;
15'b0000101010001001010 : color = 12'he73;
15'b0000101010001001011 : color = 12'he73;
15'b0000101010001001100 : color = 12'he73;
15'b0000101010001001101 : color = 12'he73;
15'b0000101010001001110 : color = 12'he73;
15'b0000101010001001111 : color = 12'he73;
15'b0000101010001010000 : color = 12'he73;
15'b0000101010001010001 : color = 12'he73;
15'b0000101010001010010 : color = 12'he73;
15'b0000101010001010011 : color = 12'he73;
15'b0000101010001010100 : color = 12'he73;
15'b0000101010001010101 : color = 12'he73;
15'b0000101010001010110 : color = 12'he73;
15'b0000101010001010111 : color = 12'he73;
15'b0000101010001011000 : color = 12'he73;
15'b0000101010001011001 : color = 12'he73;
15'b0000101010001011010 : color = 12'he73;
15'b0000101010001011011 : color = 12'he73;
15'b0000101010001011100 : color = 12'he73;
15'b0000101010001011101 : color = 12'he73;
15'b0000101010001011110 : color = 12'he73;
15'b0000101010001011111 : color = 12'he73;
15'b0000101010001100000 : color = 12'he73;
15'b0000101010001100001 : color = 12'he73;
15'b0000101010001100010 : color = 12'he73;
15'b0000101010001100011 : color = 12'he73;
15'b0000101010001100100 : color = 12'he73;
15'b0000101010001100101 : color = 12'he73;
15'b0000101010001100110 : color = 12'he73;
15'b0000101010001100111 : color = 12'he73;
15'b0000101010001101000 : color = 12'he73;
15'b0000101010001101001 : color = 12'he73;
15'b0000101010001101010 : color = 12'he73;
15'b0000101010001101011 : color = 12'he73;
15'b0000101010001101100 : color = 12'he73;
15'b0000101010001101101 : color = 12'he73;
15'b0000101010001101110 : color = 12'he73;
15'b0000101010001101111 : color = 12'he73;
15'b0000101010001110000 : color = 12'he73;
15'b0000101010001110001 : color = 12'he73;
15'b0000101010001110010 : color = 12'he73;
15'b0000101010001110011 : color = 12'he73;
15'b0000101010001110100 : color = 12'he73;
15'b0000101010001110101 : color = 12'he73;
15'b0000101010001110110 : color = 12'he73;
15'b0000101010001110111 : color = 12'he73;
15'b0000101010001111000 : color = 12'he73;
15'b0000101010001111001 : color = 12'he73;
15'b0000101010001111010 : color = 12'he73;
15'b0000101010001111011 : color = 12'he73;
15'b0000101010001111100 : color = 12'he73;
15'b0000101010001111101 : color = 12'he73;
15'b0000101010001111110 : color = 12'he73;
15'b0000101010001111111 : color = 12'he73;
15'b0000101010010000000 : color = 12'he73;
15'b0000101010010000001 : color = 12'he73;
15'b0000101010010000010 : color = 12'he73;
15'b0000101010010000011 : color = 12'he73;
15'b0000101010010000100 : color = 12'he73;
15'b0000101010010000101 : color = 12'he73;
15'b0000101010010000110 : color = 12'he73;
15'b0000101010010000111 : color = 12'he73;
15'b0000101010010001000 : color = 12'he73;
15'b0000101010010001001 : color = 12'he73;
15'b0000101010010001010 : color = 12'he73;
15'b0000101010010001011 : color = 12'he73;
15'b0000101010010001100 : color = 12'he73;
15'b0000101010010001101 : color = 12'he73;
15'b0000101010010001110 : color = 12'he73;
15'b0000101010010001111 : color = 12'he73;
15'b0000101010010010000 : color = 12'he73;
15'b0000101010010010001 : color = 12'he73;
15'b0000101010010010010 : color = 12'he73;
15'b0000101010010010011 : color = 12'he73;
15'b0000101010010010100 : color = 12'he73;
15'b0000101010010010101 : color = 12'he73;
15'b0000101010010010110 : color = 12'he73;
15'b0000101010010010111 : color = 12'he73;
15'b0000101010010011000 : color = 12'he73;
15'b0000101010010011001 : color = 12'he73;
15'b0000101010010011010 : color = 12'he73;
15'b0000101010010011011 : color = 12'he73;
15'b0000101010010011100 : color = 12'he73;
15'b0000101010010011101 : color = 12'he73;
15'b0000101010010011110 : color = 12'he73;
15'b0000101010010011111 : color = 12'he73;
15'b0000101010010100000 : color = 12'he73;
15'b0000101010010100001 : color = 12'he73;
15'b0000101010010100010 : color = 12'he73;
15'b0000101010010100011 : color = 12'he73;
15'b0000101010010100100 : color = 12'he73;
15'b0000101010010100101 : color = 12'he73;
15'b0000101010010100110 : color = 12'he73;
15'b0000101010010100111 : color = 12'he73;
15'b0000101010010101000 : color = 12'he73;
15'b0000101010010101001 : color = 12'he73;
15'b0000101010010101010 : color = 12'he73;
15'b0000101010010101011 : color = 12'he73;
15'b0000101010010101100 : color = 12'he73;
15'b0000101010010101101 : color = 12'he73;
15'b0000101010010101110 : color = 12'he73;
15'b0000101010010101111 : color = 12'he73;
15'b0000101010010110000 : color = 12'he73;
15'b0000101010010110001 : color = 12'he73;
15'b0000101010010110010 : color = 12'he73;
15'b0000101010010110011 : color = 12'he73;
15'b0000101010010110100 : color = 12'he73;
15'b0000101010010110101 : color = 12'he73;
15'b0000101010010110110 : color = 12'he73;
15'b0000101010010110111 : color = 12'he73;
15'b0000101010010111000 : color = 12'he73;
15'b0000101010010111001 : color = 12'he73;
15'b0000101010010111010 : color = 12'he73;
15'b0000101010010111011 : color = 12'he73;
15'b0000101010010111100 : color = 12'he73;
15'b0000101010010111101 : color = 12'he73;
15'b0000101010010111110 : color = 12'he73;
15'b0000101010010111111 : color = 12'he73;
15'b0000101010011000000 : color = 12'he73;
15'b0000101010011000001 : color = 12'he73;
15'b0000101010011000010 : color = 12'he73;
15'b0000101010011000011 : color = 12'he73;
15'b0000101010011000100 : color = 12'he73;
15'b0000101010011000101 : color = 12'he73;
15'b0000101010011000110 : color = 12'he73;
15'b0000101010011000111 : color = 12'he73;
15'b0000101010011001000 : color = 12'he73;
15'b0000101010011001001 : color = 12'he73;
15'b0000101010011001010 : color = 12'he73;
15'b0000101010011001011 : color = 12'he73;
15'b0000101010011001100 : color = 12'he73;
15'b0000101010011001101 : color = 12'he73;
15'b0000101010011001110 : color = 12'he73;
15'b0000101010011001111 : color = 12'he73;
15'b0000101010011010000 : color = 12'he73;
15'b0000101010011010001 : color = 12'he73;
15'b0000101010011010010 : color = 12'he73;
15'b0000101010011010011 : color = 12'he73;
15'b0000101010011010100 : color = 12'he73;
15'b0000101010011010101 : color = 12'he73;
15'b0000101010011010110 : color = 12'he73;
15'b0000101010011010111 : color = 12'he73;
15'b0000101010011011000 : color = 12'he73;
15'b0000101010011011001 : color = 12'he73;
15'b0000101010011011010 : color = 12'he73;
15'b0000101010011011011 : color = 12'he73;
15'b0000101010011011100 : color = 12'he73;
15'b0000101010011011101 : color = 12'he73;
15'b0000101010011011110 : color = 12'he73;
15'b0000101010011011111 : color = 12'he73;
15'b0000101010011100000 : color = 12'he73;
15'b0000101010011100001 : color = 12'he73;
15'b0000101010011100010 : color = 12'he73;
15'b0000101010011100011 : color = 12'he73;
15'b0000101010011100100 : color = 12'he73;
15'b0000101010011100101 : color = 12'he73;
15'b0000101010011100110 : color = 12'he73;
15'b0000101010011100111 : color = 12'he73;
15'b0000101010011101000 : color = 12'he73;
15'b0000101010011101001 : color = 12'he73;
15'b0000101010011101010 : color = 12'he73;
15'b0000101010011101011 : color = 12'he73;
15'b0000101010011101100 : color = 12'he73;
15'b0000101010011101101 : color = 12'he73;
15'b0000101010011101110 : color = 12'he73;
15'b0000101010011101111 : color = 12'he73;
15'b0000101010011110000 : color = 12'he73;
15'b0000101010011110001 : color = 12'he73;
15'b0000101010011110010 : color = 12'he73;
15'b0000101010011110011 : color = 12'he73;
15'b0000101010011110100 : color = 12'he73;
15'b0000101010011110101 : color = 12'he73;
15'b0000101010011110110 : color = 12'he73;
15'b0000101010011110111 : color = 12'he73;
15'b0000101010011111000 : color = 12'he73;
15'b0000101010011111001 : color = 12'he73;
15'b0000101010011111010 : color = 12'he73;
15'b0000101010011111011 : color = 12'he73;
15'b0000101010011111100 : color = 12'he73;
15'b0000101010011111101 : color = 12'he73;
15'b0000101010011111110 : color = 12'he73;
15'b0000101010011111111 : color = 12'he73;
15'b0000101010100000000 : color = 12'he73;
15'b0000101010100000001 : color = 12'he73;
15'b0000101010100000010 : color = 12'he73;
15'b0000101010100000011 : color = 12'he73;
15'b0000101010100000100 : color = 12'he73;
15'b0000101010100000101 : color = 12'he73;
15'b0000101010100000110 : color = 12'he73;
15'b0000101010100000111 : color = 12'he73;
15'b0000101010100001000 : color = 12'he73;
15'b0000101010100001001 : color = 12'he73;
15'b0000101010100001010 : color = 12'he73;
15'b0000101010100001011 : color = 12'he73;
15'b0000101010100001100 : color = 12'he73;
15'b0000101010100001101 : color = 12'he73;
15'b0000101010100001110 : color = 12'he73;
15'b0000101010100001111 : color = 12'he73;
15'b0000101010100010000 : color = 12'he73;
15'b0000101010100010001 : color = 12'he73;
15'b0000101010100010010 : color = 12'he73;
15'b0000101010100010011 : color = 12'he73;
15'b0000101010100010100 : color = 12'he73;
15'b0000101010100010101 : color = 12'he73;
15'b0000101010100010110 : color = 12'he73;
15'b0000101010100010111 : color = 12'he73;
15'b0000101010100011000 : color = 12'he73;
15'b0000101010100011001 : color = 12'he73;
15'b0000101010100011010 : color = 12'he73;
15'b0000101010100011011 : color = 12'he73;
15'b0000101010100011100 : color = 12'he73;
15'b0000101010100011101 : color = 12'he73;
15'b0000101010100011110 : color = 12'he73;
15'b0000101010100011111 : color = 12'he73;
15'b0000101010100100000 : color = 12'he73;
15'b0000101010100100001 : color = 12'he73;
15'b0000101010100100010 : color = 12'he73;
15'b0000101010100100011 : color = 12'he73;
15'b0000101010100100100 : color = 12'he73;
15'b0000101010100100101 : color = 12'he73;
15'b0000101010100100110 : color = 12'he73;
15'b0000101010100100111 : color = 12'he73;
15'b0000101010100101000 : color = 12'he73;
15'b0000101010100101001 : color = 12'he73;
15'b0000101010100101010 : color = 12'he73;
15'b0000101010100101011 : color = 12'he73;
15'b0000101010100101100 : color = 12'he73;
15'b0000101010100101101 : color = 12'he73;
15'b0000101010100101110 : color = 12'he73;
15'b0000101010100101111 : color = 12'he73;
15'b0000101010100110000 : color = 12'he73;
15'b0000101010100110001 : color = 12'he73;
15'b0000101010100110010 : color = 12'he73;
15'b0000101010100110011 : color = 12'he73;
15'b0000101010100110100 : color = 12'he73;
15'b0000101010100110101 : color = 12'he73;
15'b0000101010100110110 : color = 12'he73;
15'b0000101010100110111 : color = 12'he73;
15'b0000101010100111000 : color = 12'he73;
15'b0000101010100111001 : color = 12'he73;
15'b0000101010100111010 : color = 12'he73;
15'b0000101010100111011 : color = 12'he73;
15'b0000101010100111100 : color = 12'he73;
15'b0000101010100111101 : color = 12'he73;
15'b0000101010100111110 : color = 12'he73;
15'b0000101010100111111 : color = 12'he73;
15'b0000101010101000000 : color = 12'he73;
15'b0000101010101000001 : color = 12'he73;
15'b0000101010101000010 : color = 12'he73;
15'b0000101010101000011 : color = 12'he73;
15'b0000101010101000100 : color = 12'he73;
15'b0000101010101000101 : color = 12'he73;
15'b0000101010101000110 : color = 12'he73;
15'b0000101010101000111 : color = 12'he73;
15'b0000101010101001000 : color = 12'he73;
15'b0000101010101001001 : color = 12'he73;
15'b0000101010101001010 : color = 12'he73;
15'b0000101010101001011 : color = 12'he73;
15'b0000101010101001100 : color = 12'he73;
15'b0000101010101001101 : color = 12'he73;
15'b0000101010101001110 : color = 12'he73;
15'b0000101010101001111 : color = 12'he73;
15'b0000101010101010000 : color = 12'he73;
15'b0000101010101010001 : color = 12'he73;
15'b0000101010101010010 : color = 12'he73;
15'b0000101010101010011 : color = 12'he73;
15'b0000101010101010100 : color = 12'he73;
15'b0000101010101010101 : color = 12'he73;
15'b0000101010101010110 : color = 12'he73;
15'b0000101010101010111 : color = 12'he73;
15'b0000101010101011000 : color = 12'he73;
15'b0000101010101011001 : color = 12'he73;
15'b0000101010101011010 : color = 12'he73;
15'b0000101010101011011 : color = 12'he73;
15'b0000101010101011100 : color = 12'he73;
15'b0000101010101011101 : color = 12'he73;
15'b0000101010101011110 : color = 12'he73;
15'b0000101010101011111 : color = 12'he73;
15'b0000101010101100000 : color = 12'he73;
15'b0000101010101100001 : color = 12'he73;
15'b0000101010101100010 : color = 12'he73;
15'b0000101010101100011 : color = 12'he73;
15'b0000101010101100100 : color = 12'he73;
15'b0000101010101100101 : color = 12'he73;
15'b0000101010101100110 : color = 12'he73;
15'b0000101010101100111 : color = 12'he73;
15'b0000101010101101000 : color = 12'he73;
15'b0000101010101101001 : color = 12'he73;
15'b0000101010101101010 : color = 12'he73;
15'b0000101010101101011 : color = 12'he73;
15'b0000101010101101100 : color = 12'he73;
15'b0000101010101101101 : color = 12'he73;
15'b0000101010101101110 : color = 12'he73;
15'b0000101010101101111 : color = 12'he73;
15'b0000101010101110000 : color = 12'he73;
15'b0000101010101110001 : color = 12'he73;
15'b0000101010101110010 : color = 12'he73;
15'b0000101010101110011 : color = 12'he73;
15'b0000101010101110100 : color = 12'he73;
15'b0000101010101110101 : color = 12'he73;
15'b0000101010101110110 : color = 12'he73;
15'b0000101010101110111 : color = 12'he73;
15'b0000101010101111000 : color = 12'he73;
15'b0000101010101111001 : color = 12'he73;
15'b0000101010101111010 : color = 12'he73;
15'b0000101010101111011 : color = 12'he73;
15'b0000101010101111100 : color = 12'he73;
15'b0000101010101111101 : color = 12'he73;
15'b0000101010101111110 : color = 12'he73;
15'b0000101010101111111 : color = 12'he73;
15'b0000101010110000000 : color = 12'he73;
15'b0000101010110000001 : color = 12'he73;
15'b0000101010110000010 : color = 12'he73;
15'b0000101010110000011 : color = 12'he73;
15'b0000101010110000100 : color = 12'he73;
15'b0000101010110000101 : color = 12'he73;
15'b0000101010110000110 : color = 12'he73;
15'b0000101010110000111 : color = 12'he73;
15'b0000101010110001000 : color = 12'he73;
15'b0000101010110001001 : color = 12'he73;
15'b0000101010110001010 : color = 12'he73;
15'b0000101010110001011 : color = 12'he73;
15'b0000101010110001100 : color = 12'he73;
15'b0000101010110001101 : color = 12'he73;
15'b0000101010110001110 : color = 12'he73;
15'b0000101010110001111 : color = 12'he73;
15'b0000101010110010000 : color = 12'he73;
15'b0000101010110010001 : color = 12'he73;
15'b0000101010110010010 : color = 12'he73;
15'b0000101010110010011 : color = 12'he73;
15'b0000101010110010100 : color = 12'he73;
15'b0000101010110010101 : color = 12'he73;
15'b0000101010110010110 : color = 12'he73;
15'b0000101010110010111 : color = 12'he73;
15'b0000101010110011000 : color = 12'he73;
15'b0000101010110011001 : color = 12'he73;
15'b0000101010110011010 : color = 12'he73;
15'b0000101010110011011 : color = 12'he73;
15'b0000101010110011100 : color = 12'he73;
15'b0000101010110011101 : color = 12'he73;
15'b0000101010110011110 : color = 12'he73;
15'b0000101010110011111 : color = 12'he73;
15'b0000101010110100000 : color = 12'he73;
15'b0000101010110100001 : color = 12'he73;
15'b0000101010110100010 : color = 12'he73;
15'b0000101010110100011 : color = 12'he73;
15'b0000101010110100100 : color = 12'he73;
15'b0000101010110100101 : color = 12'he73;
15'b0000101010110100110 : color = 12'he73;
15'b0000101010110100111 : color = 12'he73;
15'b0000101010110101000 : color = 12'he73;
15'b0000101010110101001 : color = 12'he73;
15'b0000101010110101010 : color = 12'he73;
15'b0000101010110101011 : color = 12'he73;
15'b0000101010110101100 : color = 12'he73;
15'b0000101010110101101 : color = 12'he73;
15'b0000101001111101100 : color = 12'he73;
15'b0000101001111101101 : color = 12'he73;
15'b0000101001111101110 : color = 12'he73;
15'b0000101001111101111 : color = 12'he73;
15'b0000101001111110000 : color = 12'he73;
15'b0000101001111110001 : color = 12'he73;
15'b0000101001111110010 : color = 12'he73;
15'b0000101001111110011 : color = 12'he73;
15'b0000101001111110100 : color = 12'he73;
15'b0000101001111110101 : color = 12'he73;
15'b0000101001111110110 : color = 12'he73;
15'b0000101001111110111 : color = 12'he73;
15'b0000101001111111000 : color = 12'he73;
15'b0000101001111111001 : color = 12'he73;
15'b0000101001111111010 : color = 12'he73;
15'b0000101001111111011 : color = 12'he73;
15'b0000101001111111100 : color = 12'he73;
15'b0000101001111111101 : color = 12'he73;
15'b0000101001111111110 : color = 12'he73;
15'b0000101001111111111 : color = 12'he73;
15'b0000101010000000000 : color = 12'he73;
15'b0000101010000000001 : color = 12'he73;
15'b0000101010000000010 : color = 12'he73;
15'b0000101010000000011 : color = 12'he73;
15'b0000101010000000100 : color = 12'he73;
15'b0000101010000000101 : color = 12'he73;
15'b0000101010000000110 : color = 12'he73;
15'b0000101010000000111 : color = 12'he73;
15'b0000101010000001000 : color = 12'he73;
15'b0000101010000001001 : color = 12'he73;
15'b0000101010000001010 : color = 12'he73;
15'b0000101010000001011 : color = 12'he73;
15'b0000101010000001100 : color = 12'he73;
15'b0000101010000001101 : color = 12'he73;
15'b0000101010000001110 : color = 12'he73;
15'b0000101010000001111 : color = 12'he73;
15'b0000101010000010000 : color = 12'he73;
15'b0000101010000010001 : color = 12'he73;
15'b0000101010000010010 : color = 12'he73;
15'b0000101010000010011 : color = 12'he73;
15'b0000101010000010100 : color = 12'he73;
15'b0000101010000010101 : color = 12'he73;
15'b0000101010000010110 : color = 12'he73;
15'b0000101010000010111 : color = 12'he73;
15'b0000101010000011000 : color = 12'he73;
15'b0000101010000011001 : color = 12'he73;
15'b0000101010000011010 : color = 12'he73;
15'b0000101010000011011 : color = 12'he73;
15'b0000101010000011100 : color = 12'he73;
15'b0000101010000011101 : color = 12'he73;
15'b0000101010000011110 : color = 12'he73;
15'b0000101010000011111 : color = 12'he73;
15'b0000101010000100000 : color = 12'he73;
15'b0000101010000100001 : color = 12'he73;
15'b0000101010000100010 : color = 12'he73;
15'b0000101010000100011 : color = 12'he73;
15'b0000101010000100100 : color = 12'he73;
15'b0000101010000100101 : color = 12'he73;
15'b0000101010000100110 : color = 12'he73;
15'b0000101010000100111 : color = 12'he73;
15'b0000101010000101000 : color = 12'he73;
15'b0000101010000101001 : color = 12'he73;
15'b0000101010000101010 : color = 12'he73;
15'b0000101010000101011 : color = 12'he73;
15'b0000101010000101100 : color = 12'he73;
15'b0000101010000101101 : color = 12'he73;
15'b0000101010000101110 : color = 12'he73;
15'b0000101010000101111 : color = 12'he73;
15'b0000101010000110000 : color = 12'he73;
15'b0000101010000110001 : color = 12'he73;
15'b0000101010000110010 : color = 12'he73;
15'b0000101010000110011 : color = 12'he73;
15'b0000101010000110100 : color = 12'he73;
15'b0000101010000110101 : color = 12'he73;
15'b0000101010000110110 : color = 12'he73;
15'b0000101010000110111 : color = 12'he73;
15'b0000101010000111000 : color = 12'he73;
15'b0000101010000111001 : color = 12'he73;
15'b0000101010000111010 : color = 12'he73;
15'b0000101010000111011 : color = 12'he73;
15'b0000101010000111100 : color = 12'he73;
15'b0000101010000111101 : color = 12'he73;
15'b0000101010000111110 : color = 12'he73;
15'b0000101010000111111 : color = 12'he73;
15'b0000101010001000000 : color = 12'he73;
15'b0000101010001000001 : color = 12'he73;
15'b0000101010001000010 : color = 12'he73;
15'b0000101010001000011 : color = 12'he73;
15'b0000101010001000100 : color = 12'he73;
15'b0000101010001000101 : color = 12'he73;
15'b0000101010001000110 : color = 12'he73;
15'b0000101010001000111 : color = 12'he73;
15'b0000101010001001000 : color = 12'he73;
15'b0000101010001001001 : color = 12'he73;
15'b0000101010001001010 : color = 12'he73;
15'b0000101010001001011 : color = 12'he73;
15'b0000101010001001100 : color = 12'he73;
15'b0000101010001001101 : color = 12'he73;
15'b0000101010001001110 : color = 12'he73;
15'b0000101010001001111 : color = 12'he73;
15'b0000101010001010000 : color = 12'he73;
15'b0000101010001010001 : color = 12'he73;
15'b0000101010001010010 : color = 12'he73;
15'b0000101010001010011 : color = 12'he73;
15'b0000101010001010100 : color = 12'he73;
15'b0000101010001010101 : color = 12'he73;
15'b0000101010001010110 : color = 12'he73;
15'b0000101010001010111 : color = 12'he73;
15'b0000101010001011000 : color = 12'he73;
15'b0000101010001011001 : color = 12'he73;
15'b0000101010001011010 : color = 12'he73;
15'b0000101010001011011 : color = 12'he73;
15'b0000101010001011100 : color = 12'he73;
15'b0000101010001011101 : color = 12'he73;
15'b0000101010001011110 : color = 12'he73;
15'b0000101010001011111 : color = 12'he73;
15'b0000101010001100000 : color = 12'he73;
15'b0000101010001100001 : color = 12'he73;
15'b0000101010001100010 : color = 12'he73;
15'b0000101010001100011 : color = 12'he73;
15'b0000101010001100100 : color = 12'he73;
15'b0000101010001100101 : color = 12'he73;
15'b0000101010001100110 : color = 12'he73;
15'b0000101010001100111 : color = 12'he73;
15'b0000101010001101000 : color = 12'he73;
15'b0000101010001101001 : color = 12'he73;
15'b0000101010001101010 : color = 12'he73;
15'b0000101010001101011 : color = 12'he73;
15'b0000101010001101100 : color = 12'he73;
15'b0000101010001101101 : color = 12'he73;
15'b0000101010001101110 : color = 12'he73;
15'b0000101010001101111 : color = 12'he73;
15'b0000101010001110000 : color = 12'he73;
15'b0000101010001110001 : color = 12'he73;
15'b0000101010001110010 : color = 12'he73;
15'b0000101010001110011 : color = 12'he73;
15'b0000101010001110100 : color = 12'he73;
15'b0000101010001110101 : color = 12'he73;
15'b0000101010001110110 : color = 12'he73;
15'b0000101010001110111 : color = 12'he73;
15'b0000101010001111000 : color = 12'he73;
15'b0000101010001111001 : color = 12'he73;
15'b0000101010001111010 : color = 12'he73;
15'b0000101010001111011 : color = 12'he73;
15'b0000101010001111100 : color = 12'he73;
15'b0000101010001111101 : color = 12'he73;
15'b0000101010001111110 : color = 12'he73;
15'b0000101010001111111 : color = 12'he73;
15'b0000101010010000000 : color = 12'he73;
15'b0000101010010000001 : color = 12'he73;
15'b0000101010010000010 : color = 12'he73;
15'b0000101010010000011 : color = 12'he73;
15'b0000101010010000100 : color = 12'he73;
15'b0000101010010000101 : color = 12'he73;
15'b0000101010010000110 : color = 12'he73;
15'b0000101010010000111 : color = 12'he73;
15'b0000101010010001000 : color = 12'he73;
15'b0000101010010001001 : color = 12'he73;
15'b0000101010010001010 : color = 12'he73;
15'b0000101010010001011 : color = 12'he73;
15'b0000101010010001100 : color = 12'he73;
15'b0000101010010001101 : color = 12'he73;
15'b0000101010010001110 : color = 12'he73;
15'b0000101010010001111 : color = 12'he73;
15'b0000101010010010000 : color = 12'he73;
15'b0000101010010010001 : color = 12'he73;
15'b0000101010010010010 : color = 12'he73;
15'b0000101010010010011 : color = 12'he73;
15'b0000101010010010100 : color = 12'he73;
15'b0000101010010010101 : color = 12'he73;
15'b0000101010010010110 : color = 12'he73;
15'b0000101010010010111 : color = 12'he73;
15'b0000101010010011000 : color = 12'he73;
15'b0000101010010011001 : color = 12'he73;
15'b0000101010010011010 : color = 12'he73;
15'b0000101010010011011 : color = 12'he73;
15'b0000101010010011100 : color = 12'he73;
15'b0000101010010011101 : color = 12'he73;
15'b0000101010010011110 : color = 12'he73;
15'b0000101010010011111 : color = 12'he73;
15'b0000101010010100000 : color = 12'he73;
15'b0000101010010100001 : color = 12'he73;
15'b0000101010010100010 : color = 12'he73;
15'b0000101010010100011 : color = 12'he73;
15'b0000101010010100100 : color = 12'he73;
15'b0000101010010100101 : color = 12'he73;
15'b0000101010010100110 : color = 12'he73;
15'b0000101010010100111 : color = 12'he73;
15'b0000101010010101000 : color = 12'he73;
15'b0000101010010101001 : color = 12'he73;
15'b0000101010010101010 : color = 12'he73;
15'b0000101010010101011 : color = 12'he73;
15'b0000101010010101100 : color = 12'he73;
15'b0000101010010101101 : color = 12'he73;
15'b0000101010010101110 : color = 12'he73;
15'b0000101010010101111 : color = 12'he73;
15'b0000101010010110000 : color = 12'he73;
15'b0000101010010110001 : color = 12'he73;
15'b0000101010010110010 : color = 12'he73;
15'b0000101010010110011 : color = 12'he73;
15'b0000101010010110100 : color = 12'he73;
15'b0000101010010110101 : color = 12'he73;
15'b0000101010010110110 : color = 12'he73;
15'b0000101010010110111 : color = 12'he73;
15'b0000101010010111000 : color = 12'he73;
15'b0000101010010111001 : color = 12'he73;
15'b0000101010010111010 : color = 12'he73;
15'b0000101010010111011 : color = 12'he73;
15'b0000101010010111100 : color = 12'he73;
15'b0000101010010111101 : color = 12'he73;
15'b0000101010010111110 : color = 12'he73;
15'b0000101010010111111 : color = 12'he73;
15'b0000101010011000000 : color = 12'he73;
15'b0000101010011000001 : color = 12'he73;
15'b0000101010011000010 : color = 12'he73;
15'b0000101010011000011 : color = 12'he73;
15'b0000101010011000100 : color = 12'he73;
15'b0000101010011000101 : color = 12'he73;
15'b0000101010011000110 : color = 12'he73;
15'b0000101010011000111 : color = 12'he73;
15'b0000101010011001000 : color = 12'he73;
15'b0000101010011001001 : color = 12'he73;
15'b0000101010011001010 : color = 12'he73;
15'b0000101010011001011 : color = 12'he73;
15'b0000101010011001100 : color = 12'he73;
15'b0000101010011001101 : color = 12'he73;
15'b0000101010011001110 : color = 12'he73;
15'b0000101010011001111 : color = 12'he73;
15'b0000101010011010000 : color = 12'he73;
15'b0000101010011010001 : color = 12'he73;
15'b0000101010011010010 : color = 12'he73;
15'b0000101010011010011 : color = 12'he73;
15'b0000101010011010100 : color = 12'he73;
15'b0000101010011010101 : color = 12'he73;
15'b0000101010011010110 : color = 12'he73;
15'b0000101010011010111 : color = 12'he73;
15'b0000101010011011000 : color = 12'he73;
15'b0000101010011011001 : color = 12'he73;
15'b0000101010011011010 : color = 12'he73;
15'b0000101010011011011 : color = 12'he73;
15'b0000101010011011100 : color = 12'he73;
15'b0000101010011011101 : color = 12'he73;
15'b0000101010011011110 : color = 12'he73;
15'b0000101010011011111 : color = 12'he73;
15'b0000101010011100000 : color = 12'he73;
15'b0000101010011100001 : color = 12'he73;
15'b0000101010011100010 : color = 12'he73;
15'b0000101010011100011 : color = 12'he73;
15'b0000101010011100100 : color = 12'he73;
15'b0000101010011100101 : color = 12'he73;
15'b0000101010011100110 : color = 12'he73;
15'b0000101010011100111 : color = 12'he73;
15'b0000101010011101000 : color = 12'he73;
15'b0000101010011101001 : color = 12'he73;
15'b0000101010011101010 : color = 12'he73;
15'b0000101010011101011 : color = 12'he73;
15'b0000101010011101100 : color = 12'he73;
15'b0000101010011101101 : color = 12'he73;
15'b0000101010011101110 : color = 12'he73;
15'b0000101010011101111 : color = 12'he73;
15'b0000101010011110000 : color = 12'he73;
15'b0000101010011110001 : color = 12'he73;
15'b0000101010011110010 : color = 12'he73;
15'b0000101010011110011 : color = 12'he73;
15'b0000101010011110100 : color = 12'he73;
15'b0000101010011110101 : color = 12'he73;
15'b0000101010011110110 : color = 12'he73;
15'b0000101010011110111 : color = 12'he73;
15'b0000101010011111000 : color = 12'he73;
15'b0000101010011111001 : color = 12'he73;
15'b0000101010011111010 : color = 12'he73;
15'b0000101010011111011 : color = 12'he73;
15'b0000101010011111100 : color = 12'he73;
15'b0000101010011111101 : color = 12'he73;
15'b0000101010011111110 : color = 12'he73;
15'b0000101010011111111 : color = 12'he73;
15'b0000101010100000000 : color = 12'he73;
15'b0000101010100000001 : color = 12'he73;
15'b0000101010100000010 : color = 12'he73;
15'b0000101010100000011 : color = 12'he73;
15'b0000101010100000100 : color = 12'he73;
15'b0000101010100000101 : color = 12'he73;
15'b0000101010100000110 : color = 12'he73;
15'b0000101010100000111 : color = 12'he73;
15'b0000101010100001000 : color = 12'he73;
15'b0000101010100001001 : color = 12'he73;
15'b0000101010100001010 : color = 12'he73;
15'b0000101010100001011 : color = 12'he73;
15'b0000101010100001100 : color = 12'he73;
15'b0000101010100001101 : color = 12'he73;
15'b0000101010100001110 : color = 12'he73;
15'b0000101010100001111 : color = 12'he73;
15'b0000101010100010000 : color = 12'he73;
15'b0000101010100010001 : color = 12'he73;
15'b0000101010100010010 : color = 12'he73;
15'b0000101010100010011 : color = 12'he73;
15'b0000101010100010100 : color = 12'he73;
15'b0000101010100010101 : color = 12'he73;
15'b0000101010100010110 : color = 12'he73;
15'b0000101010100010111 : color = 12'he73;
15'b0000101010100011000 : color = 12'he73;
15'b0000101010100011001 : color = 12'he73;
15'b0000101010100011010 : color = 12'he73;
15'b0000101010100011011 : color = 12'he73;
15'b0000101010100011100 : color = 12'he73;
15'b0000101010100011101 : color = 12'he73;
15'b0000101010100011110 : color = 12'he73;
15'b0000101010100011111 : color = 12'he73;
15'b0000101010100100000 : color = 12'he73;
15'b0000101010100100001 : color = 12'he73;
15'b0000101010100100010 : color = 12'he73;
15'b0000101010100100011 : color = 12'he73;
15'b0000101010100100100 : color = 12'he73;
15'b0000101010100100101 : color = 12'he73;
15'b0000101010100100110 : color = 12'he73;
15'b0000101010100100111 : color = 12'he73;
15'b0000101010100101000 : color = 12'he73;
15'b0000101010100101001 : color = 12'he73;
15'b0000101010100101010 : color = 12'he73;
15'b0000101010100101011 : color = 12'he73;
15'b0000101010100101100 : color = 12'he73;
15'b0000101010100101101 : color = 12'he73;
15'b0000101010100101110 : color = 12'he73;
15'b0000101010100101111 : color = 12'he73;
15'b0000101010100110000 : color = 12'he73;
15'b0000101010100110001 : color = 12'he73;
15'b0000101010100110010 : color = 12'he73;
15'b0000101010100110011 : color = 12'he73;
15'b0000101010100110100 : color = 12'he73;
15'b0000101010100110101 : color = 12'he73;
15'b0000101010100110110 : color = 12'he73;
15'b0000101010100110111 : color = 12'he73;
15'b0000101010100111000 : color = 12'he73;
15'b0000101010100111001 : color = 12'he73;
15'b0000101010100111010 : color = 12'he73;
15'b0000101010100111011 : color = 12'he73;
15'b0000101010100111100 : color = 12'he73;
15'b0000101010100111101 : color = 12'he73;
15'b0000101010100111110 : color = 12'he73;
15'b0000101010100111111 : color = 12'he73;
15'b0000101010101000000 : color = 12'he73;
15'b0000101010101000001 : color = 12'he73;
15'b0000101010101000010 : color = 12'he73;
15'b0000101010101000011 : color = 12'he73;
15'b0000101010101000100 : color = 12'he73;
15'b0000101010101000101 : color = 12'he73;
15'b0000101010101000110 : color = 12'he73;
15'b0000101010101000111 : color = 12'he73;
15'b0000101010101001000 : color = 12'he73;
15'b0000101010101001001 : color = 12'he73;
15'b0000101010101001010 : color = 12'he73;
15'b0000101010101001011 : color = 12'he73;
15'b0000101010101001100 : color = 12'he73;
15'b0000101010101001101 : color = 12'he73;
15'b0000101010101001110 : color = 12'he73;
15'b0000101010101001111 : color = 12'he73;
15'b0000101010101010000 : color = 12'he73;
15'b0000101010101010001 : color = 12'he73;
15'b0000101010101010010 : color = 12'he73;
15'b0000101010101010011 : color = 12'he73;
15'b0000101010101010100 : color = 12'he73;
15'b0000101010101010101 : color = 12'he73;
15'b0000101010101010110 : color = 12'he73;
15'b0000101010101010111 : color = 12'he73;
15'b0000101010101011000 : color = 12'he73;
15'b0000101010101011001 : color = 12'he73;
15'b0000101010101011010 : color = 12'he73;
15'b0000101010101011011 : color = 12'he73;
15'b0000101010101011100 : color = 12'he73;
15'b0000101010101011101 : color = 12'he73;
15'b0000101010101011110 : color = 12'he73;
15'b0000101010101011111 : color = 12'he73;
15'b0000101010101100000 : color = 12'he73;
15'b0000101010101100001 : color = 12'he73;
15'b0000101010101100010 : color = 12'he73;
15'b0000101010101100011 : color = 12'he73;
15'b0000101010101100100 : color = 12'he73;
15'b0000101010101100101 : color = 12'he73;
15'b0000101010101100110 : color = 12'he73;
15'b0000101010101100111 : color = 12'he73;
15'b0000101010101101000 : color = 12'he73;
15'b0000101010101101001 : color = 12'he73;
15'b0000101010101101010 : color = 12'he73;
15'b0000101010101101011 : color = 12'he73;
15'b0000101010101101100 : color = 12'he73;
15'b0000101010101101101 : color = 12'he73;
15'b0000101010101101110 : color = 12'he73;
15'b0000101010101101111 : color = 12'he73;
15'b0000101010101110000 : color = 12'he73;
15'b0000101010101110001 : color = 12'he73;
15'b0000101010101110010 : color = 12'he73;
15'b0000101010101110011 : color = 12'he73;
15'b0000101010101110100 : color = 12'he73;
15'b0000101010101110101 : color = 12'he73;
15'b0000101010101110110 : color = 12'he73;
15'b0000101010101110111 : color = 12'he73;
15'b0000101010101111000 : color = 12'he73;
15'b0000101010101111001 : color = 12'he73;
15'b0000101010101111010 : color = 12'he73;
15'b0000101010101111011 : color = 12'he73;
15'b0000101010101111100 : color = 12'he73;
15'b0000101010101111101 : color = 12'he73;
15'b0000101010101111110 : color = 12'he73;
15'b0000101010101111111 : color = 12'he73;
15'b0000101010110000000 : color = 12'he73;
15'b0000101010110000001 : color = 12'he73;
15'b0000101010110000010 : color = 12'he73;
15'b0000101010110000011 : color = 12'he73;
15'b0000101010110000100 : color = 12'he73;
15'b0000101010110000101 : color = 12'he73;
15'b0000101010110000110 : color = 12'he73;
15'b0000101010110000111 : color = 12'he73;
15'b0000101010110001000 : color = 12'he73;
15'b0000101010110001001 : color = 12'he73;
15'b0000101010110001010 : color = 12'he73;
15'b0000101010110001011 : color = 12'he73;
15'b0000101010110001100 : color = 12'he73;
15'b0000101010110001101 : color = 12'he73;
15'b0000101010110001110 : color = 12'he73;
15'b0000101010110001111 : color = 12'he73;
15'b0000101010110010000 : color = 12'he73;
15'b0000101010110010001 : color = 12'he73;
15'b0000101010110010010 : color = 12'he73;
15'b0000101010110010011 : color = 12'he73;
15'b0000101010110010100 : color = 12'he73;
15'b0000101010110010101 : color = 12'he73;
15'b0000101010110010110 : color = 12'he73;
15'b0000101010110010111 : color = 12'he73;
15'b0000101010110011000 : color = 12'he73;
15'b0000101010110011001 : color = 12'he73;
15'b0000101010110011010 : color = 12'he73;
15'b0000101010110011011 : color = 12'he73;
15'b0000101010110011100 : color = 12'he73;
15'b0000101010110011101 : color = 12'he73;
15'b0000101010110011110 : color = 12'he73;
15'b0000101010110011111 : color = 12'he73;
15'b0000101010110100000 : color = 12'he73;
15'b0000101010110100001 : color = 12'he73;
15'b0000101010110100010 : color = 12'he73;
15'b0000101010110100011 : color = 12'he73;
15'b0000101010110100100 : color = 12'he73;
15'b0000101010110100101 : color = 12'he73;
15'b0000101010110100110 : color = 12'he73;
15'b0000101010110100111 : color = 12'he73;
15'b0000101010110101000 : color = 12'he73;
15'b0000101010110101001 : color = 12'he73;
15'b0000101010110101010 : color = 12'he73;
15'b0000101010110101011 : color = 12'he73;
15'b0000101010110101100 : color = 12'he73;
15'b0000101010110101101 : color = 12'he73;
15'b0000101010110101110 : color = 12'he73;
15'b0000101010110101111 : color = 12'he73;
15'b0000101010110110000 : color = 12'he73;
15'b0000101010110110001 : color = 12'he73;
15'b0000101010110110010 : color = 12'he73;
15'b0000101010110110011 : color = 12'he73;
15'b0000101010110110100 : color = 12'he73;
15'b0000101010110110101 : color = 12'he73;
15'b0000101010110110110 : color = 12'he73;
15'b0000101010110110111 : color = 12'he73;
15'b0000101010110111000 : color = 12'he73;
15'b0000101010110111001 : color = 12'he73;
15'b0000101010110111010 : color = 12'he73;
15'b0000101010110111011 : color = 12'he73;
15'b0000101010110111100 : color = 12'he73;
15'b0000101010110111101 : color = 12'he73;
15'b0000101010110111110 : color = 12'he73;
15'b0000101010110111111 : color = 12'he73;
15'b0000101010111000000 : color = 12'he73;
15'b0000101010111000001 : color = 12'he73;
15'b0000101010111000010 : color = 12'he73;
15'b0000101010111000011 : color = 12'he73;
15'b0000101010111000100 : color = 12'he73;
15'b0000101010111000101 : color = 12'he73;
15'b0000101010111000110 : color = 12'he73;
15'b0000101010111000111 : color = 12'he73;
15'b0000101010111001000 : color = 12'he73;
15'b0000101010111001001 : color = 12'he73;
15'b0000101010111001010 : color = 12'he73;
15'b0000101010111001011 : color = 12'he73;
15'b0000101010111001100 : color = 12'he73;
15'b0000101010111001101 : color = 12'he73;
15'b0000101010111001110 : color = 12'he73;
15'b0000101010111001111 : color = 12'he73;
15'b0000101010111010000 : color = 12'he73;
15'b0000101010111010001 : color = 12'he73;
15'b0000101010111010010 : color = 12'he73;
15'b0000101010111010011 : color = 12'he73;
15'b0000101010111010100 : color = 12'he73;
15'b0000101010111010101 : color = 12'he73;
15'b0000101010111010110 : color = 12'he73;
15'b0000101010000010101 : color = 12'he73;
15'b0000101010000010110 : color = 12'he73;
15'b0000101010000010111 : color = 12'he73;
15'b0000101010000011000 : color = 12'he73;
15'b0000101010000011001 : color = 12'he73;
15'b0000101010000011010 : color = 12'he73;
15'b0000101010000011011 : color = 12'he73;
15'b0000101010000011100 : color = 12'he73;
15'b0000101010000011101 : color = 12'he73;
15'b0000101010000011110 : color = 12'he73;
15'b0000101010000011111 : color = 12'he73;
15'b0000101010000100000 : color = 12'he73;
15'b0000101010000100001 : color = 12'he73;
15'b0000101010000100010 : color = 12'he73;
15'b0000101010000100011 : color = 12'he73;
15'b0000101010000100100 : color = 12'he73;
15'b0000101010000100101 : color = 12'he73;
15'b0000101010000100110 : color = 12'he73;
15'b0000101010000100111 : color = 12'he73;
15'b0000101010000101000 : color = 12'he73;
15'b0000101010000101001 : color = 12'he73;
15'b0000101010000101010 : color = 12'he73;
15'b0000101010000101011 : color = 12'he73;
15'b0000101010000101100 : color = 12'he73;
15'b0000101010000101101 : color = 12'he73;
15'b0000101010000101110 : color = 12'he73;
15'b0000101010000101111 : color = 12'he73;
15'b0000101010000110000 : color = 12'he73;
15'b0000101010000110001 : color = 12'he73;
15'b0000101010000110010 : color = 12'he73;
15'b0000101010000110011 : color = 12'he73;
15'b0000101010000110100 : color = 12'he73;
15'b0000101010000110101 : color = 12'he73;
15'b0000101010000110110 : color = 12'he73;
15'b0000101010000110111 : color = 12'he73;
15'b0000101010000111000 : color = 12'he73;
15'b0000101010000111001 : color = 12'he73;
15'b0000101010000111010 : color = 12'he73;
15'b0000101010000111011 : color = 12'he73;
15'b0000101010000111100 : color = 12'he73;
15'b0000101010000111101 : color = 12'he73;
15'b0000101010000111110 : color = 12'he73;
15'b0000101010000111111 : color = 12'he73;
15'b0000101010001000000 : color = 12'he73;
15'b0000101010001000001 : color = 12'he73;
15'b0000101010001000010 : color = 12'he73;
15'b0000101010001000011 : color = 12'he73;
15'b0000101010001000100 : color = 12'he73;
15'b0000101010001000101 : color = 12'he73;
15'b0000101010001000110 : color = 12'he73;
15'b0000101010001000111 : color = 12'he73;
15'b0000101010001001000 : color = 12'he73;
15'b0000101010001001001 : color = 12'he73;
15'b0000101010001001010 : color = 12'he73;
15'b0000101010001001011 : color = 12'he73;
15'b0000101010001001100 : color = 12'he73;
15'b0000101010001001101 : color = 12'he73;
15'b0000101010001001110 : color = 12'he73;
15'b0000101010001001111 : color = 12'he73;
15'b0000101010001010000 : color = 12'he73;
15'b0000101010001010001 : color = 12'he73;
15'b0000101010001010010 : color = 12'he73;
15'b0000101010001010011 : color = 12'he73;
15'b0000101010001010100 : color = 12'he73;
15'b0000101010001010101 : color = 12'he73;
15'b0000101010001010110 : color = 12'he73;
15'b0000101010001010111 : color = 12'he73;
15'b0000101010001011000 : color = 12'he73;
15'b0000101010001011001 : color = 12'he73;
15'b0000101010001011010 : color = 12'he73;
15'b0000101010001011011 : color = 12'he73;
15'b0000101010001011100 : color = 12'he73;
15'b0000101010001011101 : color = 12'he73;
15'b0000101010001011110 : color = 12'he73;
15'b0000101010001011111 : color = 12'he73;
15'b0000101010001100000 : color = 12'he73;
15'b0000101010001100001 : color = 12'he73;
15'b0000101010001100010 : color = 12'he73;
15'b0000101010001100011 : color = 12'he73;
15'b0000101010001100100 : color = 12'he73;
15'b0000101010001100101 : color = 12'he73;
15'b0000101010001100110 : color = 12'he73;
15'b0000101010001100111 : color = 12'he73;
15'b0000101010001101000 : color = 12'he73;
15'b0000101010001101001 : color = 12'he73;
15'b0000101010001101010 : color = 12'he73;
15'b0000101010001101011 : color = 12'he73;
15'b0000101010001101100 : color = 12'he73;
15'b0000101010001101101 : color = 12'he73;
15'b0000101010001101110 : color = 12'he73;
15'b0000101010001101111 : color = 12'he73;
15'b0000101010001110000 : color = 12'he73;
15'b0000101010001110001 : color = 12'he73;
15'b0000101010001110010 : color = 12'he73;
15'b0000101010001110011 : color = 12'he73;
15'b0000101010001110100 : color = 12'he73;
15'b0000101010001110101 : color = 12'he73;
15'b0000101010001110110 : color = 12'he73;
15'b0000101010001110111 : color = 12'he73;
15'b0000101010001111000 : color = 12'he73;
15'b0000101010001111001 : color = 12'he73;
15'b0000101010001111010 : color = 12'he73;
15'b0000101010001111011 : color = 12'he73;
15'b0000101010001111100 : color = 12'he73;
15'b0000101010001111101 : color = 12'he73;
15'b0000101010001111110 : color = 12'he73;
15'b0000101010001111111 : color = 12'he73;
15'b0000101010010000000 : color = 12'he73;
15'b0000101010010000001 : color = 12'he73;
15'b0000101010010000010 : color = 12'he73;
15'b0000101010010000011 : color = 12'he73;
15'b0000101010010000100 : color = 12'he73;
15'b0000101010010000101 : color = 12'he73;
15'b0000101010010000110 : color = 12'he73;
15'b0000101010010000111 : color = 12'he73;
15'b0000101010010001000 : color = 12'he73;
15'b0000101010010001001 : color = 12'he73;
15'b0000101010010001010 : color = 12'he73;
15'b0000101010010001011 : color = 12'he73;
15'b0000101010010001100 : color = 12'he73;
15'b0000101010010001101 : color = 12'he73;
15'b0000101010010001110 : color = 12'he73;
15'b0000101010010001111 : color = 12'he73;
15'b0000101010010010000 : color = 12'he73;
15'b0000101010010010001 : color = 12'he73;
15'b0000101010010010010 : color = 12'he73;
15'b0000101010010010011 : color = 12'he73;
15'b0000101010010010100 : color = 12'he73;
15'b0000101010010010101 : color = 12'he73;
15'b0000101010010010110 : color = 12'he73;
15'b0000101010010010111 : color = 12'he73;
15'b0000101010010011000 : color = 12'he73;
15'b0000101010010011001 : color = 12'he73;
15'b0000101010010011010 : color = 12'he73;
15'b0000101010010011011 : color = 12'he73;
15'b0000101010010011100 : color = 12'he73;
15'b0000101010010011101 : color = 12'he73;
15'b0000101010010011110 : color = 12'he73;
15'b0000101010010011111 : color = 12'he73;
15'b0000101010010100000 : color = 12'he73;
15'b0000101010010100001 : color = 12'he73;
15'b0000101010010100010 : color = 12'he73;
15'b0000101010010100011 : color = 12'he73;
15'b0000101010010100100 : color = 12'he73;
15'b0000101010010100101 : color = 12'he73;
15'b0000101010010100110 : color = 12'he73;
15'b0000101010010100111 : color = 12'he73;
15'b0000101010010101000 : color = 12'he73;
15'b0000101010010101001 : color = 12'he73;
15'b0000101010010101010 : color = 12'he73;
15'b0000101010010101011 : color = 12'he73;
15'b0000101010010101100 : color = 12'he73;
15'b0000101010010101101 : color = 12'he73;
15'b0000101010010101110 : color = 12'he73;
15'b0000101010010101111 : color = 12'he73;
15'b0000101010010110000 : color = 12'he73;
15'b0000101010010110001 : color = 12'he73;
15'b0000101010010110010 : color = 12'he73;
15'b0000101010010110011 : color = 12'he73;
15'b0000101010010110100 : color = 12'he73;
15'b0000101010010110101 : color = 12'he73;
15'b0000101010010110110 : color = 12'he73;
15'b0000101010010110111 : color = 12'he73;
15'b0000101010010111000 : color = 12'he73;
15'b0000101010010111001 : color = 12'he73;
15'b0000101010010111010 : color = 12'he73;
15'b0000101010010111011 : color = 12'he73;
15'b0000101010010111100 : color = 12'he73;
15'b0000101010010111101 : color = 12'he73;
15'b0000101010010111110 : color = 12'he73;
15'b0000101010010111111 : color = 12'he73;
15'b0000101010011000000 : color = 12'he73;
15'b0000101010011000001 : color = 12'he73;
15'b0000101010011000010 : color = 12'he73;
15'b0000101010011000011 : color = 12'he73;
15'b0000101010011000100 : color = 12'he73;
15'b0000101010011000101 : color = 12'he73;
15'b0000101010011000110 : color = 12'he73;
15'b0000101010011000111 : color = 12'he73;
15'b0000101010011001000 : color = 12'he73;
15'b0000101010011001001 : color = 12'he73;
15'b0000101010011001010 : color = 12'he73;
15'b0000101010011001011 : color = 12'he73;
15'b0000101010011001100 : color = 12'he73;
15'b0000101010011001101 : color = 12'he73;
15'b0000101010011001110 : color = 12'he73;
15'b0000101010011001111 : color = 12'he73;
15'b0000101010011010000 : color = 12'he73;
15'b0000101010011010001 : color = 12'he73;
15'b0000101010011010010 : color = 12'he73;
15'b0000101010011010011 : color = 12'he73;
15'b0000101010011010100 : color = 12'he73;
15'b0000101010011010101 : color = 12'he73;
15'b0000101010011010110 : color = 12'he73;
15'b0000101010011010111 : color = 12'he73;
15'b0000101010011011000 : color = 12'he73;
15'b0000101010011011001 : color = 12'he73;
15'b0000101010011011010 : color = 12'he73;
15'b0000101010011011011 : color = 12'he73;
15'b0000101010011011100 : color = 12'he73;
15'b0000101010011011101 : color = 12'he73;
15'b0000101010011011110 : color = 12'he73;
15'b0000101010011011111 : color = 12'he73;
15'b0000101010011100000 : color = 12'he73;
15'b0000101010011100001 : color = 12'he73;
15'b0000101010011100010 : color = 12'he73;
15'b0000101010011100011 : color = 12'he73;
15'b0000101010011100100 : color = 12'he73;
15'b0000101010011100101 : color = 12'he73;
15'b0000101010011100110 : color = 12'he73;
15'b0000101010011100111 : color = 12'he73;
15'b0000101010011101000 : color = 12'he73;
15'b0000101010011101001 : color = 12'he73;
15'b0000101010011101010 : color = 12'he73;
15'b0000101010011101011 : color = 12'he73;
15'b0000101010011101100 : color = 12'he73;
15'b0000101010011101101 : color = 12'he73;
15'b0000101010011101110 : color = 12'he73;
15'b0000101010011101111 : color = 12'he73;
15'b0000101010011110000 : color = 12'he73;
15'b0000101010011110001 : color = 12'he73;
15'b0000101010011110010 : color = 12'he73;
15'b0000101010011110011 : color = 12'he73;
15'b0000101010011110100 : color = 12'he73;
15'b0000101010011110101 : color = 12'he73;
15'b0000101010011110110 : color = 12'he73;
15'b0000101010011110111 : color = 12'he73;
15'b0000101010011111000 : color = 12'he73;
15'b0000101010011111001 : color = 12'he73;
15'b0000101010011111010 : color = 12'he73;
15'b0000101010011111011 : color = 12'he73;
15'b0000101010011111100 : color = 12'he73;
15'b0000101010011111101 : color = 12'he73;
15'b0000101010011111110 : color = 12'he73;
15'b0000101010011111111 : color = 12'he73;
15'b0000101010100000000 : color = 12'he73;
15'b0000101010100000001 : color = 12'he73;
15'b0000101010100000010 : color = 12'he73;
15'b0000101010100000011 : color = 12'he73;
15'b0000101010100000100 : color = 12'he73;
15'b0000101010100000101 : color = 12'he73;
15'b0000101010100000110 : color = 12'he73;
15'b0000101010100000111 : color = 12'he73;
15'b0000101010100001000 : color = 12'he73;
15'b0000101010100001001 : color = 12'he73;
15'b0000101010100001010 : color = 12'he73;
15'b0000101010100001011 : color = 12'he73;
15'b0000101010100001100 : color = 12'he73;
15'b0000101010100001101 : color = 12'he73;
15'b0000101010100001110 : color = 12'he73;
15'b0000101010100001111 : color = 12'he73;
15'b0000101010100010000 : color = 12'he73;
15'b0000101010100010001 : color = 12'he73;
15'b0000101010100010010 : color = 12'he73;
15'b0000101010100010011 : color = 12'he73;
15'b0000101010100010100 : color = 12'he73;
15'b0000101010100010101 : color = 12'he73;
15'b0000101010100010110 : color = 12'he73;
15'b0000101010100010111 : color = 12'he73;
15'b0000101010100011000 : color = 12'he73;
15'b0000101010100011001 : color = 12'he73;
15'b0000101010100011010 : color = 12'he73;
15'b0000101010100011011 : color = 12'he73;
15'b0000101010100011100 : color = 12'he73;
15'b0000101010100011101 : color = 12'he73;
15'b0000101010100011110 : color = 12'he73;
15'b0000101010100011111 : color = 12'he73;
15'b0000101010100100000 : color = 12'he73;
15'b0000101010100100001 : color = 12'he73;
15'b0000101010100100010 : color = 12'he73;
15'b0000101010100100011 : color = 12'he73;
15'b0000101010100100100 : color = 12'he73;
15'b0000101010100100101 : color = 12'he73;
15'b0000101010100100110 : color = 12'he73;
15'b0000101010100100111 : color = 12'he73;
15'b0000101010100101000 : color = 12'he73;
15'b0000101010100101001 : color = 12'he73;
15'b0000101010100101010 : color = 12'he73;
15'b0000101010100101011 : color = 12'he73;
15'b0000101010100101100 : color = 12'he73;
15'b0000101010100101101 : color = 12'he73;
15'b0000101010100101110 : color = 12'he73;
15'b0000101010100101111 : color = 12'he73;
15'b0000101010100110000 : color = 12'he73;
15'b0000101010100110001 : color = 12'he73;
15'b0000101010100110010 : color = 12'he73;
15'b0000101010100110011 : color = 12'he73;
15'b0000101010100110100 : color = 12'he73;
15'b0000101010100110101 : color = 12'he73;
15'b0000101010100110110 : color = 12'he73;
15'b0000101010100110111 : color = 12'he73;
15'b0000101010100111000 : color = 12'he73;
15'b0000101010100111001 : color = 12'he73;
15'b0000101010100111010 : color = 12'he73;
15'b0000101010100111011 : color = 12'he73;
15'b0000101010100111100 : color = 12'he73;
15'b0000101010100111101 : color = 12'he73;
15'b0000101010100111110 : color = 12'he73;
15'b0000101010100111111 : color = 12'he73;
15'b0000101010101000000 : color = 12'he73;
15'b0000101010101000001 : color = 12'he73;
15'b0000101010101000010 : color = 12'he73;
15'b0000101010101000011 : color = 12'he73;
15'b0000101010101000100 : color = 12'he73;
15'b0000101010101000101 : color = 12'he73;
15'b0000101010101000110 : color = 12'he73;
15'b0000101010101000111 : color = 12'he73;
15'b0000101010101001000 : color = 12'he73;
15'b0000101010101001001 : color = 12'he73;
15'b0000101010101001010 : color = 12'he73;
15'b0000101010101001011 : color = 12'he73;
15'b0000101010101001100 : color = 12'he73;
15'b0000101010101001101 : color = 12'he73;
15'b0000101010101001110 : color = 12'he73;
15'b0000101010101001111 : color = 12'he73;
15'b0000101010101010000 : color = 12'he73;
15'b0000101010101010001 : color = 12'he73;
15'b0000101010101010010 : color = 12'he73;
15'b0000101010101010011 : color = 12'he73;
15'b0000101010101010100 : color = 12'he73;
15'b0000101010101010101 : color = 12'he73;
15'b0000101010101010110 : color = 12'he73;
15'b0000101010101010111 : color = 12'he73;
15'b0000101010101011000 : color = 12'he73;
15'b0000101010101011001 : color = 12'he73;
15'b0000101010101011010 : color = 12'he73;
15'b0000101010101011011 : color = 12'he73;
15'b0000101010101011100 : color = 12'he73;
15'b0000101010101011101 : color = 12'he73;
15'b0000101010101011110 : color = 12'he73;
15'b0000101010101011111 : color = 12'he73;
15'b0000101010101100000 : color = 12'he73;
15'b0000101010101100001 : color = 12'he73;
15'b0000101010101100010 : color = 12'he73;
15'b0000101010101100011 : color = 12'he73;
15'b0000101010101100100 : color = 12'he73;
15'b0000101010101100101 : color = 12'he73;
15'b0000101010101100110 : color = 12'he73;
15'b0000101010101100111 : color = 12'he73;
15'b0000101010101101000 : color = 12'he73;
15'b0000101010101101001 : color = 12'he73;
15'b0000101010101101010 : color = 12'he73;
15'b0000101010101101011 : color = 12'he73;
15'b0000101010101101100 : color = 12'he73;
15'b0000101010101101101 : color = 12'he73;
15'b0000101010101101110 : color = 12'he73;
15'b0000101010101101111 : color = 12'he73;
15'b0000101010101110000 : color = 12'he73;
15'b0000101010101110001 : color = 12'he73;
15'b0000101010101110010 : color = 12'he73;
15'b0000101010101110011 : color = 12'he73;
15'b0000101010101110100 : color = 12'he73;
15'b0000101010101110101 : color = 12'he73;
15'b0000101010101110110 : color = 12'he73;
15'b0000101010101110111 : color = 12'he73;
15'b0000101010101111000 : color = 12'he73;
15'b0000101010101111001 : color = 12'he73;
15'b0000101010101111010 : color = 12'he73;
15'b0000101010101111011 : color = 12'he73;
15'b0000101010101111100 : color = 12'he73;
15'b0000101010101111101 : color = 12'he73;
15'b0000101010101111110 : color = 12'he73;
15'b0000101010101111111 : color = 12'he73;
15'b0000101010110000000 : color = 12'he73;
15'b0000101010110000001 : color = 12'he73;
15'b0000101010110000010 : color = 12'he73;
15'b0000101010110000011 : color = 12'he73;
15'b0000101010110000100 : color = 12'he73;
15'b0000101010110000101 : color = 12'he73;
15'b0000101010110000110 : color = 12'he73;
15'b0000101010110000111 : color = 12'he73;
15'b0000101010110001000 : color = 12'he73;
15'b0000101010110001001 : color = 12'he73;
15'b0000101010110001010 : color = 12'he73;
15'b0000101010110001011 : color = 12'he73;
15'b0000101010110001100 : color = 12'he73;
15'b0000101010110001101 : color = 12'he73;
15'b0000101010110001110 : color = 12'he73;
15'b0000101010110001111 : color = 12'he73;
15'b0000101010110010000 : color = 12'he73;
15'b0000101010110010001 : color = 12'he73;
15'b0000101010110010010 : color = 12'he73;
15'b0000101010110010011 : color = 12'he73;
15'b0000101010110010100 : color = 12'he73;
15'b0000101010110010101 : color = 12'he73;
15'b0000101010110010110 : color = 12'he73;
15'b0000101010110010111 : color = 12'he73;
15'b0000101010110011000 : color = 12'he73;
15'b0000101010110011001 : color = 12'he73;
15'b0000101010110011010 : color = 12'he73;
15'b0000101010110011011 : color = 12'he73;
15'b0000101010110011100 : color = 12'he73;
15'b0000101010110011101 : color = 12'he73;
15'b0000101010110011110 : color = 12'he73;
15'b0000101010110011111 : color = 12'he73;
15'b0000101010110100000 : color = 12'he73;
15'b0000101010110100001 : color = 12'he73;
15'b0000101010110100010 : color = 12'he73;
15'b0000101010110100011 : color = 12'he73;
15'b0000101010110100100 : color = 12'he73;
15'b0000101010110100101 : color = 12'he73;
15'b0000101010110100110 : color = 12'he73;
15'b0000101010110100111 : color = 12'he73;
15'b0000101010110101000 : color = 12'he73;
15'b0000101010110101001 : color = 12'he73;
15'b0000101010110101010 : color = 12'he73;
15'b0000101010110101011 : color = 12'he73;
15'b0000101010110101100 : color = 12'he73;
15'b0000101010110101101 : color = 12'he73;
15'b0000101010110101110 : color = 12'he73;
15'b0000101010110101111 : color = 12'he73;
15'b0000101010110110000 : color = 12'he73;
15'b0000101010110110001 : color = 12'he73;
15'b0000101010110110010 : color = 12'he73;
15'b0000101010110110011 : color = 12'he73;
15'b0000101010110110100 : color = 12'he73;
15'b0000101010110110101 : color = 12'he73;
15'b0000101010110110110 : color = 12'he73;
15'b0000101010110110111 : color = 12'he73;
15'b0000101010110111000 : color = 12'he73;
15'b0000101010110111001 : color = 12'he73;
15'b0000101010110111010 : color = 12'he73;
15'b0000101010110111011 : color = 12'he73;
15'b0000101010110111100 : color = 12'he73;
15'b0000101010110111101 : color = 12'he73;
15'b0000101010110111110 : color = 12'he73;
15'b0000101010110111111 : color = 12'he73;
15'b0000101010111000000 : color = 12'he73;
15'b0000101010111000001 : color = 12'he73;
15'b0000101010111000010 : color = 12'he73;
15'b0000101010111000011 : color = 12'he73;
15'b0000101010111000100 : color = 12'he73;
15'b0000101010111000101 : color = 12'he73;
15'b0000101010111000110 : color = 12'he73;
15'b0000101010111000111 : color = 12'he73;
15'b0000101010111001000 : color = 12'he73;
15'b0000101010111001001 : color = 12'he73;
15'b0000101010111001010 : color = 12'he73;
15'b0000101010111001011 : color = 12'he73;
15'b0000101010111001100 : color = 12'he73;
15'b0000101010111001101 : color = 12'he73;
15'b0000101010111001110 : color = 12'he73;
15'b0000101010111001111 : color = 12'he73;
15'b0000101010111010000 : color = 12'he73;
15'b0000101010111010001 : color = 12'he73;
15'b0000101010111010010 : color = 12'he73;
15'b0000101010111010011 : color = 12'he73;
15'b0000101010111010100 : color = 12'he73;
15'b0000101010111010101 : color = 12'he73;
15'b0000101010111010110 : color = 12'he73;
15'b0000101010111010111 : color = 12'he73;
15'b0000101010111011000 : color = 12'he73;
15'b0000101010111011001 : color = 12'he73;
15'b0000101010111011010 : color = 12'he73;
15'b0000101010111011011 : color = 12'he73;
15'b0000101010111011100 : color = 12'he73;
15'b0000101010111011101 : color = 12'he73;
15'b0000101010111011110 : color = 12'he73;
15'b0000101010111011111 : color = 12'he73;
15'b0000101010111100000 : color = 12'he73;
15'b0000101010111100001 : color = 12'he73;
15'b0000101010111100010 : color = 12'he73;
15'b0000101010111100011 : color = 12'he73;
15'b0000101010111100100 : color = 12'he73;
15'b0000101010111100101 : color = 12'he73;
15'b0000101010111100110 : color = 12'he73;
15'b0000101010111100111 : color = 12'he73;
15'b0000101010111101000 : color = 12'he73;
15'b0000101010111101001 : color = 12'he73;
15'b0000101010111101010 : color = 12'he73;
15'b0000101010111101011 : color = 12'he73;
15'b0000101010111101100 : color = 12'he73;
15'b0000101010111101101 : color = 12'he73;
15'b0000101010111101110 : color = 12'he73;
15'b0000101010111101111 : color = 12'he73;
15'b0000101010111110000 : color = 12'he73;
15'b0000101010111110001 : color = 12'he73;
15'b0000101010111110010 : color = 12'he73;
15'b0000101010111110011 : color = 12'he73;
15'b0000101010111110100 : color = 12'he73;
15'b0000101010111110101 : color = 12'he73;
15'b0000101010111110110 : color = 12'he73;
15'b0000101010111110111 : color = 12'he73;
15'b0000101010111111000 : color = 12'he73;
15'b0000101010111111001 : color = 12'he73;
15'b0000101010111111010 : color = 12'he73;
15'b0000101010111111011 : color = 12'he73;
15'b0000101010111111100 : color = 12'he73;
15'b0000101010111111101 : color = 12'he73;
15'b0000101010111111110 : color = 12'he73;
15'b0000101010111111111 : color = 12'he73;
15'b0000101010000111110 : color = 12'he73;
15'b0000101010000111111 : color = 12'he73;
15'b0000101010001000000 : color = 12'he73;
15'b0000101010001000001 : color = 12'he73;
15'b0000101010001000010 : color = 12'he73;
15'b0000101010001000011 : color = 12'he73;
15'b0000101010001000100 : color = 12'he73;
15'b0000101010001000101 : color = 12'he73;
15'b0000101010001000110 : color = 12'he73;
15'b0000101010001000111 : color = 12'he73;
15'b0000101010001001000 : color = 12'he73;
15'b0000101010001001001 : color = 12'he73;
15'b0000101010001001010 : color = 12'he73;
15'b0000101010001001011 : color = 12'he73;
15'b0000101010001001100 : color = 12'he73;
15'b0000101010001001101 : color = 12'he73;
15'b0000101010001001110 : color = 12'he73;
15'b0000101010001001111 : color = 12'he73;
15'b0000101010001010000 : color = 12'he73;
15'b0000101010001010001 : color = 12'he73;
15'b0000101010001010010 : color = 12'he73;
15'b0000101010001010011 : color = 12'he73;
15'b0000101010001010100 : color = 12'he73;
15'b0000101010001010101 : color = 12'he73;
15'b0000101010001010110 : color = 12'he73;
15'b0000101010001010111 : color = 12'he73;
15'b0000101010001011000 : color = 12'he73;
15'b0000101010001011001 : color = 12'he73;
15'b0000101010001011010 : color = 12'he73;
15'b0000101010001011011 : color = 12'he73;
15'b0000101010001011100 : color = 12'he73;
15'b0000101010001011101 : color = 12'he73;
15'b0000101010001011110 : color = 12'he73;
15'b0000101010001011111 : color = 12'he73;
15'b0000101010001100000 : color = 12'he73;
15'b0000101010001100001 : color = 12'he73;
15'b0000101010001100010 : color = 12'he73;
15'b0000101010001100011 : color = 12'he73;
15'b0000101010001100100 : color = 12'he73;
15'b0000101010001100101 : color = 12'he73;
15'b0000101010001100110 : color = 12'he73;
15'b0000101010001100111 : color = 12'he73;
15'b0000101010001101000 : color = 12'he73;
15'b0000101010001101001 : color = 12'he73;
15'b0000101010001101010 : color = 12'he73;
15'b0000101010001101011 : color = 12'he73;
15'b0000101010001101100 : color = 12'he73;
15'b0000101010001101101 : color = 12'he73;
15'b0000101010001101110 : color = 12'he73;
15'b0000101010001101111 : color = 12'he73;
15'b0000101010001110000 : color = 12'he73;
15'b0000101010001110001 : color = 12'he73;
15'b0000101010001110010 : color = 12'he73;
15'b0000101010001110011 : color = 12'he73;
15'b0000101010001110100 : color = 12'he73;
15'b0000101010001110101 : color = 12'he73;
15'b0000101010001110110 : color = 12'he73;
15'b0000101010001110111 : color = 12'he73;
15'b0000101010001111000 : color = 12'he73;
15'b0000101010001111001 : color = 12'he73;
15'b0000101010001111010 : color = 12'he73;
15'b0000101010001111011 : color = 12'he73;
15'b0000101010001111100 : color = 12'he73;
15'b0000101010001111101 : color = 12'he73;
15'b0000101010001111110 : color = 12'he73;
15'b0000101010001111111 : color = 12'he73;
15'b0000101010010000000 : color = 12'he73;
15'b0000101010010000001 : color = 12'he73;
15'b0000101010010000010 : color = 12'he73;
15'b0000101010010000011 : color = 12'he73;
15'b0000101010010000100 : color = 12'he73;
15'b0000101010010000101 : color = 12'he73;
15'b0000101010010000110 : color = 12'he73;
15'b0000101010010000111 : color = 12'he73;
15'b0000101010010001000 : color = 12'he73;
15'b0000101010010001001 : color = 12'he73;
15'b0000101010010001010 : color = 12'he73;
15'b0000101010010001011 : color = 12'he73;
15'b0000101010010001100 : color = 12'he73;
15'b0000101010010001101 : color = 12'he73;
15'b0000101010010001110 : color = 12'he73;
15'b0000101010010001111 : color = 12'he73;
15'b0000101010010010000 : color = 12'he73;
15'b0000101010010010001 : color = 12'he73;
15'b0000101010010010010 : color = 12'he73;
15'b0000101010010010011 : color = 12'he73;
15'b0000101010010010100 : color = 12'he73;
15'b0000101010010010101 : color = 12'he73;
15'b0000101010010010110 : color = 12'he73;
15'b0000101010010010111 : color = 12'he73;
15'b0000101010010011000 : color = 12'he73;
15'b0000101010010011001 : color = 12'he73;
15'b0000101010010011010 : color = 12'he73;
15'b0000101010010011011 : color = 12'he73;
15'b0000101010010011100 : color = 12'he73;
15'b0000101010010011101 : color = 12'he73;
15'b0000101010010011110 : color = 12'he73;
15'b0000101010010011111 : color = 12'he73;
15'b0000101010010100000 : color = 12'he73;
15'b0000101010010100001 : color = 12'he73;
15'b0000101010010100010 : color = 12'he73;
15'b0000101010010100011 : color = 12'he73;
15'b0000101010010100100 : color = 12'he73;
15'b0000101010010100101 : color = 12'he73;
15'b0000101010010100110 : color = 12'he73;
15'b0000101010010100111 : color = 12'he73;
15'b0000101010010101000 : color = 12'he73;
15'b0000101010010101001 : color = 12'he73;
15'b0000101010010101010 : color = 12'he73;
15'b0000101010010101011 : color = 12'he73;
15'b0000101010010101100 : color = 12'he73;
15'b0000101010010101101 : color = 12'he73;
15'b0000101010010101110 : color = 12'he73;
15'b0000101010010101111 : color = 12'he73;
15'b0000101010010110000 : color = 12'he73;
15'b0000101010010110001 : color = 12'he73;
15'b0000101010010110010 : color = 12'he73;
15'b0000101010010110011 : color = 12'he73;
15'b0000101010010110100 : color = 12'he73;
15'b0000101010010110101 : color = 12'he73;
15'b0000101010010110110 : color = 12'he73;
15'b0000101010010110111 : color = 12'he73;
15'b0000101010010111000 : color = 12'he73;
15'b0000101010010111001 : color = 12'he73;
15'b0000101010010111010 : color = 12'he73;
15'b0000101010010111011 : color = 12'he73;
15'b0000101010010111100 : color = 12'he73;
15'b0000101010010111101 : color = 12'he73;
15'b0000101010010111110 : color = 12'he73;
15'b0000101010010111111 : color = 12'he73;
15'b0000101010011000000 : color = 12'he73;
15'b0000101010011000001 : color = 12'he73;
15'b0000101010011000010 : color = 12'he73;
15'b0000101010011000011 : color = 12'he73;
15'b0000101010011000100 : color = 12'he73;
15'b0000101010011000101 : color = 12'he73;
15'b0000101010011000110 : color = 12'he73;
15'b0000101010011000111 : color = 12'he73;
15'b0000101010011001000 : color = 12'he73;
15'b0000101010011001001 : color = 12'he73;
15'b0000101010011001010 : color = 12'he73;
15'b0000101010011001011 : color = 12'he73;
15'b0000101010011001100 : color = 12'he73;
15'b0000101010011001101 : color = 12'he73;
15'b0000101010011001110 : color = 12'he73;
15'b0000101010011001111 : color = 12'he73;
15'b0000101010011010000 : color = 12'he73;
15'b0000101010011010001 : color = 12'he73;
15'b0000101010011010010 : color = 12'he73;
15'b0000101010011010011 : color = 12'he73;
15'b0000101010011010100 : color = 12'he73;
15'b0000101010011010101 : color = 12'he73;
15'b0000101010011010110 : color = 12'he73;
15'b0000101010011010111 : color = 12'he73;
15'b0000101010011011000 : color = 12'he73;
15'b0000101010011011001 : color = 12'he73;
15'b0000101010011011010 : color = 12'he73;
15'b0000101010011011011 : color = 12'he73;
15'b0000101010011011100 : color = 12'he73;
15'b0000101010011011101 : color = 12'he73;
15'b0000101010011011110 : color = 12'he73;
15'b0000101010011011111 : color = 12'he73;
15'b0000101010011100000 : color = 12'he73;
15'b0000101010011100001 : color = 12'he73;
15'b0000101010011100010 : color = 12'he73;
15'b0000101010011100011 : color = 12'he73;
15'b0000101010011100100 : color = 12'he73;
15'b0000101010011100101 : color = 12'he73;
15'b0000101010011100110 : color = 12'he73;
15'b0000101010011100111 : color = 12'he73;
15'b0000101010011101000 : color = 12'he73;
15'b0000101010011101001 : color = 12'he73;
15'b0000101010011101010 : color = 12'he73;
15'b0000101010011101011 : color = 12'he73;
15'b0000101010011101100 : color = 12'he73;
15'b0000101010011101101 : color = 12'he73;
15'b0000101010011101110 : color = 12'he73;
15'b0000101010011101111 : color = 12'he73;
15'b0000101010011110000 : color = 12'he73;
15'b0000101010011110001 : color = 12'he73;
15'b0000101010011110010 : color = 12'he73;
15'b0000101010011110011 : color = 12'he73;
15'b0000101010011110100 : color = 12'he73;
15'b0000101010011110101 : color = 12'he73;
15'b0000101010011110110 : color = 12'he73;
15'b0000101010011110111 : color = 12'he73;
15'b0000101010011111000 : color = 12'he73;
15'b0000101010011111001 : color = 12'he73;
15'b0000101010011111010 : color = 12'he73;
15'b0000101010011111011 : color = 12'he73;
15'b0000101010011111100 : color = 12'he73;
15'b0000101010011111101 : color = 12'he73;
15'b0000101010011111110 : color = 12'he73;
15'b0000101010011111111 : color = 12'he73;
15'b0000101010100000000 : color = 12'he73;
15'b0000101010100000001 : color = 12'he73;
15'b0000101010100000010 : color = 12'he73;
15'b0000101010100000011 : color = 12'he73;
15'b0000101010100000100 : color = 12'he73;
15'b0000101010100000101 : color = 12'he73;
15'b0000101010100000110 : color = 12'he73;
15'b0000101010100000111 : color = 12'he73;
15'b0000101010100001000 : color = 12'he73;
15'b0000101010100001001 : color = 12'he73;
15'b0000101010100001010 : color = 12'he73;
15'b0000101010100001011 : color = 12'he73;
15'b0000101010100001100 : color = 12'he73;
15'b0000101010100001101 : color = 12'he73;
15'b0000101010100001110 : color = 12'he73;
15'b0000101010100001111 : color = 12'he73;
15'b0000101010100010000 : color = 12'he73;
15'b0000101010100010001 : color = 12'he73;
15'b0000101010100010010 : color = 12'he73;
15'b0000101010100010011 : color = 12'he73;
15'b0000101010100010100 : color = 12'he73;
15'b0000101010100010101 : color = 12'he73;
15'b0000101010100010110 : color = 12'he73;
15'b0000101010100010111 : color = 12'he73;
15'b0000101010100011000 : color = 12'he73;
15'b0000101010100011001 : color = 12'he73;
15'b0000101010100011010 : color = 12'he73;
15'b0000101010100011011 : color = 12'he73;
15'b0000101010100011100 : color = 12'he73;
15'b0000101010100011101 : color = 12'he73;
15'b0000101010100011110 : color = 12'he73;
15'b0000101010100011111 : color = 12'he73;
15'b0000101010100100000 : color = 12'he73;
15'b0000101010100100001 : color = 12'he73;
15'b0000101010100100010 : color = 12'he73;
15'b0000101010100100011 : color = 12'he73;
15'b0000101010100100100 : color = 12'he73;
15'b0000101010100100101 : color = 12'he73;
15'b0000101010100100110 : color = 12'he73;
15'b0000101010100100111 : color = 12'he73;
15'b0000101010100101000 : color = 12'he73;
15'b0000101010100101001 : color = 12'he73;
15'b0000101010100101010 : color = 12'he73;
15'b0000101010100101011 : color = 12'he73;
15'b0000101010100101100 : color = 12'he73;
15'b0000101010100101101 : color = 12'he73;
15'b0000101010100101110 : color = 12'he73;
15'b0000101010100101111 : color = 12'he73;
15'b0000101010100110000 : color = 12'he73;
15'b0000101010100110001 : color = 12'he73;
15'b0000101010100110010 : color = 12'he73;
15'b0000101010100110011 : color = 12'he73;
15'b0000101010100110100 : color = 12'he73;
15'b0000101010100110101 : color = 12'he73;
15'b0000101010100110110 : color = 12'he73;
15'b0000101010100110111 : color = 12'he73;
15'b0000101010100111000 : color = 12'he73;
15'b0000101010100111001 : color = 12'he73;
15'b0000101010100111010 : color = 12'he73;
15'b0000101010100111011 : color = 12'he73;
15'b0000101010100111100 : color = 12'he73;
15'b0000101010100111101 : color = 12'he73;
15'b0000101010100111110 : color = 12'he73;
15'b0000101010100111111 : color = 12'he73;
15'b0000101010101000000 : color = 12'he73;
15'b0000101010101000001 : color = 12'he73;
15'b0000101010101000010 : color = 12'he73;
15'b0000101010101000011 : color = 12'he73;
15'b0000101010101000100 : color = 12'he73;
15'b0000101010101000101 : color = 12'he73;
15'b0000101010101000110 : color = 12'he73;
15'b0000101010101000111 : color = 12'he73;
15'b0000101010101001000 : color = 12'he73;
15'b0000101010101001001 : color = 12'he73;
15'b0000101010101001010 : color = 12'he73;
15'b0000101010101001011 : color = 12'he73;
15'b0000101010101001100 : color = 12'he73;
15'b0000101010101001101 : color = 12'he73;
15'b0000101010101001110 : color = 12'he73;
15'b0000101010101001111 : color = 12'he73;
15'b0000101010101010000 : color = 12'he73;
15'b0000101010101010001 : color = 12'he73;
15'b0000101010101010010 : color = 12'he73;
15'b0000101010101010011 : color = 12'he73;
15'b0000101010101010100 : color = 12'he73;
15'b0000101010101010101 : color = 12'he73;
15'b0000101010101010110 : color = 12'he73;
15'b0000101010101010111 : color = 12'he73;
15'b0000101010101011000 : color = 12'he73;
15'b0000101010101011001 : color = 12'he73;
15'b0000101010101011010 : color = 12'he73;
15'b0000101010101011011 : color = 12'he73;
15'b0000101010101011100 : color = 12'he73;
15'b0000101010101011101 : color = 12'he73;
15'b0000101010101011110 : color = 12'he73;
15'b0000101010101011111 : color = 12'he73;
15'b0000101010101100000 : color = 12'he73;
15'b0000101010101100001 : color = 12'he73;
15'b0000101010101100010 : color = 12'he73;
15'b0000101010101100011 : color = 12'he73;
15'b0000101010101100100 : color = 12'he73;
15'b0000101010101100101 : color = 12'he73;
15'b0000101010101100110 : color = 12'he73;
15'b0000101010101100111 : color = 12'he73;
15'b0000101010101101000 : color = 12'he73;
15'b0000101010101101001 : color = 12'he73;
15'b0000101010101101010 : color = 12'he73;
15'b0000101010101101011 : color = 12'he73;
15'b0000101010101101100 : color = 12'he73;
15'b0000101010101101101 : color = 12'he73;
15'b0000101010101101110 : color = 12'he73;
15'b0000101010101101111 : color = 12'he73;
15'b0000101010101110000 : color = 12'he73;
15'b0000101010101110001 : color = 12'he73;
15'b0000101010101110010 : color = 12'he73;
15'b0000101010101110011 : color = 12'he73;
15'b0000101010101110100 : color = 12'he73;
15'b0000101010101110101 : color = 12'he73;
15'b0000101010101110110 : color = 12'he73;
15'b0000101010101110111 : color = 12'he73;
15'b0000101010101111000 : color = 12'he73;
15'b0000101010101111001 : color = 12'he73;
15'b0000101010101111010 : color = 12'he73;
15'b0000101010101111011 : color = 12'he73;
15'b0000101010101111100 : color = 12'he73;
15'b0000101010101111101 : color = 12'he73;
15'b0000101010101111110 : color = 12'he73;
15'b0000101010101111111 : color = 12'he73;
15'b0000101010110000000 : color = 12'he73;
15'b0000101010110000001 : color = 12'he73;
15'b0000101010110000010 : color = 12'he73;
15'b0000101010110000011 : color = 12'he73;
15'b0000101010110000100 : color = 12'he73;
15'b0000101010110000101 : color = 12'he73;
15'b0000101010110000110 : color = 12'he73;
15'b0000101010110000111 : color = 12'he73;
15'b0000101010110001000 : color = 12'he73;
15'b0000101010110001001 : color = 12'he73;
15'b0000101010110001010 : color = 12'he73;
15'b0000101010110001011 : color = 12'he73;
15'b0000101010110001100 : color = 12'he73;
15'b0000101010110001101 : color = 12'he73;
15'b0000101010110001110 : color = 12'he73;
15'b0000101010110001111 : color = 12'he73;
15'b0000101010110010000 : color = 12'he73;
15'b0000101010110010001 : color = 12'he73;
15'b0000101010110010010 : color = 12'he73;
15'b0000101010110010011 : color = 12'he73;
15'b0000101010110010100 : color = 12'he73;
15'b0000101010110010101 : color = 12'he73;
15'b0000101010110010110 : color = 12'he73;
15'b0000101010110010111 : color = 12'he73;
15'b0000101010110011000 : color = 12'he73;
15'b0000101010110011001 : color = 12'he73;
15'b0000101010110011010 : color = 12'he73;
15'b0000101010110011011 : color = 12'he73;
15'b0000101010110011100 : color = 12'he73;
15'b0000101010110011101 : color = 12'he73;
15'b0000101010110011110 : color = 12'he73;
15'b0000101010110011111 : color = 12'he73;
15'b0000101010110100000 : color = 12'he73;
15'b0000101010110100001 : color = 12'he73;
15'b0000101010110100010 : color = 12'he73;
15'b0000101010110100011 : color = 12'he73;
15'b0000101010110100100 : color = 12'he73;
15'b0000101010110100101 : color = 12'he73;
15'b0000101010110100110 : color = 12'he73;
15'b0000101010110100111 : color = 12'he73;
15'b0000101010110101000 : color = 12'he73;
15'b0000101010110101001 : color = 12'he73;
15'b0000101010110101010 : color = 12'he73;
15'b0000101010110101011 : color = 12'he73;
15'b0000101010110101100 : color = 12'he73;
15'b0000101010110101101 : color = 12'he73;
15'b0000101010110101110 : color = 12'he73;
15'b0000101010110101111 : color = 12'he73;
15'b0000101010110110000 : color = 12'he73;
15'b0000101010110110001 : color = 12'he73;
15'b0000101010110110010 : color = 12'he73;
15'b0000101010110110011 : color = 12'he73;
15'b0000101010110110100 : color = 12'he73;
15'b0000101010110110101 : color = 12'he73;
15'b0000101010110110110 : color = 12'he73;
15'b0000101010110110111 : color = 12'he73;
15'b0000101010110111000 : color = 12'he73;
15'b0000101010110111001 : color = 12'he73;
15'b0000101010110111010 : color = 12'he73;
15'b0000101010110111011 : color = 12'he73;
15'b0000101010110111100 : color = 12'he73;
15'b0000101010110111101 : color = 12'he73;
15'b0000101010110111110 : color = 12'he73;
15'b0000101010110111111 : color = 12'he73;
15'b0000101010111000000 : color = 12'he73;
15'b0000101010111000001 : color = 12'he73;
15'b0000101010111000010 : color = 12'he73;
15'b0000101010111000011 : color = 12'he73;
15'b0000101010111000100 : color = 12'he73;
15'b0000101010111000101 : color = 12'he73;
15'b0000101010111000110 : color = 12'he73;
15'b0000101010111000111 : color = 12'he73;
15'b0000101010111001000 : color = 12'he73;
15'b0000101010111001001 : color = 12'he73;
15'b0000101010111001010 : color = 12'he73;
15'b0000101010111001011 : color = 12'he73;
15'b0000101010111001100 : color = 12'he73;
15'b0000101010111001101 : color = 12'he73;
15'b0000101010111001110 : color = 12'he73;
15'b0000101010111001111 : color = 12'he73;
15'b0000101010111010000 : color = 12'he73;
15'b0000101010111010001 : color = 12'he73;
15'b0000101010111010010 : color = 12'he73;
15'b0000101010111010011 : color = 12'he73;
15'b0000101010111010100 : color = 12'he73;
15'b0000101010111010101 : color = 12'he73;
15'b0000101010111010110 : color = 12'he73;
15'b0000101010111010111 : color = 12'he73;
15'b0000101010111011000 : color = 12'he73;
15'b0000101010111011001 : color = 12'he73;
15'b0000101010111011010 : color = 12'he73;
15'b0000101010111011011 : color = 12'he73;
15'b0000101010111011100 : color = 12'he73;
15'b0000101010111011101 : color = 12'he73;
15'b0000101010111011110 : color = 12'he73;
15'b0000101010111011111 : color = 12'he73;
15'b0000101010111100000 : color = 12'he73;
15'b0000101010111100001 : color = 12'he73;
15'b0000101010111100010 : color = 12'he73;
15'b0000101010111100011 : color = 12'he73;
15'b0000101010111100100 : color = 12'he73;
15'b0000101010111100101 : color = 12'he73;
15'b0000101010111100110 : color = 12'he73;
15'b0000101010111100111 : color = 12'he73;
15'b0000101010111101000 : color = 12'he73;
15'b0000101010111101001 : color = 12'he73;
15'b0000101010111101010 : color = 12'he73;
15'b0000101010111101011 : color = 12'he73;
15'b0000101010111101100 : color = 12'he73;
15'b0000101010111101101 : color = 12'he73;
15'b0000101010111101110 : color = 12'he73;
15'b0000101010111101111 : color = 12'he73;
15'b0000101010111110000 : color = 12'he73;
15'b0000101010111110001 : color = 12'he73;
15'b0000101010111110010 : color = 12'he73;
15'b0000101010111110011 : color = 12'he73;
15'b0000101010111110100 : color = 12'he73;
15'b0000101010111110101 : color = 12'he73;
15'b0000101010111110110 : color = 12'he73;
15'b0000101010111110111 : color = 12'he73;
15'b0000101010111111000 : color = 12'he73;
15'b0000101010111111001 : color = 12'he73;
15'b0000101010111111010 : color = 12'he73;
15'b0000101010111111011 : color = 12'he73;
15'b0000101010111111100 : color = 12'he73;
15'b0000101010111111101 : color = 12'he73;
15'b0000101010111111110 : color = 12'he73;
15'b0000101010111111111 : color = 12'he73;
15'b0000101011000000000 : color = 12'he73;
15'b0000101011000000001 : color = 12'he73;
15'b0000101011000000010 : color = 12'he73;
15'b0000101011000000011 : color = 12'he73;
15'b0000101011000000100 : color = 12'he73;
15'b0000101011000000101 : color = 12'he73;
15'b0000101011000000110 : color = 12'he73;
15'b0000101011000000111 : color = 12'he73;
15'b0000101011000001000 : color = 12'he73;
15'b0000101011000001001 : color = 12'he73;
15'b0000101011000001010 : color = 12'he73;
15'b0000101011000001011 : color = 12'he73;
15'b0000101011000001100 : color = 12'he73;
15'b0000101011000001101 : color = 12'he73;
15'b0000101011000001110 : color = 12'he73;
15'b0000101011000001111 : color = 12'he73;
15'b0000101011000010000 : color = 12'he73;
15'b0000101011000010001 : color = 12'he73;
15'b0000101011000010010 : color = 12'he73;
15'b0000101011000010011 : color = 12'he73;
15'b0000101011000010100 : color = 12'he73;
15'b0000101011000010101 : color = 12'he73;
15'b0000101011000010110 : color = 12'he73;
15'b0000101011000010111 : color = 12'he73;
15'b0000101011000011000 : color = 12'he73;
15'b0000101011000011001 : color = 12'he73;
15'b0000101011000011010 : color = 12'he73;
15'b0000101011000011011 : color = 12'he73;
15'b0000101011000011100 : color = 12'he73;
15'b0000101011000011101 : color = 12'he73;
15'b0000101011000011110 : color = 12'he73;
15'b0000101011000011111 : color = 12'he73;
15'b0000101011000100000 : color = 12'he73;
15'b0000101011000100001 : color = 12'he73;
15'b0000101011000100010 : color = 12'he73;
15'b0000101011000100011 : color = 12'he73;
15'b0000101011000100100 : color = 12'he73;
15'b0000101011000100101 : color = 12'he73;
15'b0000101011000100110 : color = 12'he73;
15'b0000101011000100111 : color = 12'he73;
15'b0000101011000101000 : color = 12'he73;
15'b0000101010001100111 : color = 12'he73;
15'b0000101010001101000 : color = 12'he73;
15'b0000101010001101001 : color = 12'he73;
15'b0000101010001101010 : color = 12'he73;
15'b0000101010001101011 : color = 12'he73;
15'b0000101010001101100 : color = 12'he73;
15'b0000101010001101101 : color = 12'he73;
15'b0000101010001101110 : color = 12'he73;
15'b0000101010001101111 : color = 12'he73;
15'b0000101010001110000 : color = 12'he73;
15'b0000101010001110001 : color = 12'he73;
15'b0000101010001110010 : color = 12'he73;
15'b0000101010001110011 : color = 12'he73;
15'b0000101010001110100 : color = 12'he73;
15'b0000101010001110101 : color = 12'he73;
15'b0000101010001110110 : color = 12'he73;
15'b0000101010001110111 : color = 12'he73;
15'b0000101010001111000 : color = 12'he73;
15'b0000101010001111001 : color = 12'he73;
15'b0000101010001111010 : color = 12'he73;
15'b0000101010001111011 : color = 12'he73;
15'b0000101010001111100 : color = 12'he73;
15'b0000101010001111101 : color = 12'he73;
15'b0000101010001111110 : color = 12'he73;
15'b0000101010001111111 : color = 12'he73;
15'b0000101010010000000 : color = 12'he73;
15'b0000101010010000001 : color = 12'he73;
15'b0000101010010000010 : color = 12'he73;
15'b0000101010010000011 : color = 12'he73;
15'b0000101010010000100 : color = 12'he73;
15'b0000101010010000101 : color = 12'he73;
15'b0000101010010000110 : color = 12'he73;
15'b0000101010010000111 : color = 12'he73;
15'b0000101010010001000 : color = 12'he73;
15'b0000101010010001001 : color = 12'he73;
15'b0000101010010001010 : color = 12'he73;
15'b0000101010010001011 : color = 12'he73;
15'b0000101010010001100 : color = 12'he73;
15'b0000101010010001101 : color = 12'he73;
15'b0000101010010001110 : color = 12'he73;
15'b0000101010010001111 : color = 12'he73;
15'b0000101010010010000 : color = 12'he73;
15'b0000101010010010001 : color = 12'he73;
15'b0000101010010010010 : color = 12'he73;
15'b0000101010010010011 : color = 12'he73;
15'b0000101010010010100 : color = 12'he73;
15'b0000101010010010101 : color = 12'he73;
15'b0000101010010010110 : color = 12'he73;
15'b0000101010010010111 : color = 12'he73;
15'b0000101010010011000 : color = 12'he73;
15'b0000101010010011001 : color = 12'he73;
15'b0000101010010011010 : color = 12'he73;
15'b0000101010010011011 : color = 12'he73;
15'b0000101010010011100 : color = 12'he73;
15'b0000101010010011101 : color = 12'he73;
15'b0000101010010011110 : color = 12'he73;
15'b0000101010010011111 : color = 12'he73;
15'b0000101010010100000 : color = 12'he73;
15'b0000101010010100001 : color = 12'he73;
15'b0000101010010100010 : color = 12'he73;
15'b0000101010010100011 : color = 12'he73;
15'b0000101010010100100 : color = 12'he73;
15'b0000101010010100101 : color = 12'he73;
15'b0000101010010100110 : color = 12'he73;
15'b0000101010010100111 : color = 12'he73;
15'b0000101010010101000 : color = 12'he73;
15'b0000101010010101001 : color = 12'he73;
15'b0000101010010101010 : color = 12'he73;
15'b0000101010010101011 : color = 12'he73;
15'b0000101010010101100 : color = 12'he73;
15'b0000101010010101101 : color = 12'he73;
15'b0000101010010101110 : color = 12'he73;
15'b0000101010010101111 : color = 12'he73;
15'b0000101010010110000 : color = 12'he73;
15'b0000101010010110001 : color = 12'he73;
15'b0000101010010110010 : color = 12'he73;
15'b0000101010010110011 : color = 12'he73;
15'b0000101010010110100 : color = 12'he73;
15'b0000101010010110101 : color = 12'he73;
15'b0000101010010110110 : color = 12'he73;
15'b0000101010010110111 : color = 12'he73;
15'b0000101010010111000 : color = 12'he73;
15'b0000101010010111001 : color = 12'he73;
15'b0000101010010111010 : color = 12'he73;
15'b0000101010010111011 : color = 12'he73;
15'b0000101010010111100 : color = 12'he73;
15'b0000101010010111101 : color = 12'he73;
15'b0000101010010111110 : color = 12'he73;
15'b0000101010010111111 : color = 12'he73;
15'b0000101010011000000 : color = 12'he73;
15'b0000101010011000001 : color = 12'he73;
15'b0000101010011000010 : color = 12'he73;
15'b0000101010011000011 : color = 12'he73;
15'b0000101010011000100 : color = 12'he73;
15'b0000101010011000101 : color = 12'he73;
15'b0000101010011000110 : color = 12'he73;
15'b0000101010011000111 : color = 12'he73;
15'b0000101010011001000 : color = 12'he73;
15'b0000101010011001001 : color = 12'he73;
15'b0000101010011001010 : color = 12'he73;
15'b0000101010011001011 : color = 12'he73;
15'b0000101010011001100 : color = 12'he73;
15'b0000101010011001101 : color = 12'he73;
15'b0000101010011001110 : color = 12'he73;
15'b0000101010011001111 : color = 12'he73;
15'b0000101010011010000 : color = 12'he73;
15'b0000101010011010001 : color = 12'he73;
15'b0000101010011010010 : color = 12'he73;
15'b0000101010011010011 : color = 12'he73;
15'b0000101010011010100 : color = 12'he73;
15'b0000101010011010101 : color = 12'he73;
15'b0000101010011010110 : color = 12'he73;
15'b0000101010011010111 : color = 12'he73;
15'b0000101010011011000 : color = 12'he73;
15'b0000101010011011001 : color = 12'he73;
15'b0000101010011011010 : color = 12'he73;
15'b0000101010011011011 : color = 12'he73;
15'b0000101010011011100 : color = 12'he73;
15'b0000101010011011101 : color = 12'he73;
15'b0000101010011011110 : color = 12'he73;
15'b0000101010011011111 : color = 12'he73;
15'b0000101010011100000 : color = 12'he73;
15'b0000101010011100001 : color = 12'he73;
15'b0000101010011100010 : color = 12'he73;
15'b0000101010011100011 : color = 12'he73;
15'b0000101010011100100 : color = 12'he73;
15'b0000101010011100101 : color = 12'he73;
15'b0000101010011100110 : color = 12'he73;
15'b0000101010011100111 : color = 12'he73;
15'b0000101010011101000 : color = 12'he73;
15'b0000101010011101001 : color = 12'he73;
15'b0000101010011101010 : color = 12'he73;
15'b0000101010011101011 : color = 12'he73;
15'b0000101010011101100 : color = 12'he73;
15'b0000101010011101101 : color = 12'he73;
15'b0000101010011101110 : color = 12'he73;
15'b0000101010011101111 : color = 12'he73;
15'b0000101010011110000 : color = 12'he73;
15'b0000101010011110001 : color = 12'he73;
15'b0000101010011110010 : color = 12'he73;
15'b0000101010011110011 : color = 12'he73;
15'b0000101010011110100 : color = 12'he73;
15'b0000101010011110101 : color = 12'he73;
15'b0000101010011110110 : color = 12'he73;
15'b0000101010011110111 : color = 12'he73;
15'b0000101010011111000 : color = 12'he73;
15'b0000101010011111001 : color = 12'he73;
15'b0000101010011111010 : color = 12'he73;
15'b0000101010011111011 : color = 12'he73;
15'b0000101010011111100 : color = 12'he73;
15'b0000101010011111101 : color = 12'he73;
15'b0000101010011111110 : color = 12'he73;
15'b0000101010011111111 : color = 12'he73;
15'b0000101010100000000 : color = 12'he73;
15'b0000101010100000001 : color = 12'he73;
15'b0000101010100000010 : color = 12'he73;
15'b0000101010100000011 : color = 12'he73;
15'b0000101010100000100 : color = 12'he73;
15'b0000101010100000101 : color = 12'he73;
15'b0000101010100000110 : color = 12'he73;
15'b0000101010100000111 : color = 12'he73;
15'b0000101010100001000 : color = 12'he73;
15'b0000101010100001001 : color = 12'he73;
15'b0000101010100001010 : color = 12'he73;
15'b0000101010100001011 : color = 12'he73;
15'b0000101010100001100 : color = 12'he73;
15'b0000101010100001101 : color = 12'he73;
15'b0000101010100001110 : color = 12'he73;
15'b0000101010100001111 : color = 12'he73;
15'b0000101010100010000 : color = 12'he73;
15'b0000101010100010001 : color = 12'he73;
15'b0000101010100010010 : color = 12'he73;
15'b0000101010100010011 : color = 12'he73;
15'b0000101010100010100 : color = 12'he73;
15'b0000101010100010101 : color = 12'he73;
15'b0000101010100010110 : color = 12'he73;
15'b0000101010100010111 : color = 12'he73;
15'b0000101010100011000 : color = 12'he73;
15'b0000101010100011001 : color = 12'he73;
15'b0000101010100011010 : color = 12'he73;
15'b0000101010100011011 : color = 12'he73;
15'b0000101010100011100 : color = 12'he73;
15'b0000101010100011101 : color = 12'he73;
15'b0000101010100011110 : color = 12'he73;
15'b0000101010100011111 : color = 12'he73;
15'b0000101010100100000 : color = 12'he73;
15'b0000101010100100001 : color = 12'he73;
15'b0000101010100100010 : color = 12'he73;
15'b0000101010100100011 : color = 12'he73;
15'b0000101010100100100 : color = 12'he73;
15'b0000101010100100101 : color = 12'he73;
15'b0000101010100100110 : color = 12'he73;
15'b0000101010100100111 : color = 12'he73;
15'b0000101010100101000 : color = 12'he73;
15'b0000101010100101001 : color = 12'he73;
15'b0000101010100101010 : color = 12'he73;
15'b0000101010100101011 : color = 12'he73;
15'b0000101010100101100 : color = 12'he73;
15'b0000101010100101101 : color = 12'he73;
15'b0000101010100101110 : color = 12'he73;
15'b0000101010100101111 : color = 12'he73;
15'b0000101010100110000 : color = 12'he73;
15'b0000101010100110001 : color = 12'he73;
15'b0000101010100110010 : color = 12'he73;
15'b0000101010100110011 : color = 12'he73;
15'b0000101010100110100 : color = 12'he73;
15'b0000101010100110101 : color = 12'he73;
15'b0000101010100110110 : color = 12'he73;
15'b0000101010100110111 : color = 12'he73;
15'b0000101010100111000 : color = 12'he73;
15'b0000101010100111001 : color = 12'he73;
15'b0000101010100111010 : color = 12'he73;
15'b0000101010100111011 : color = 12'he73;
15'b0000101010100111100 : color = 12'he73;
15'b0000101010100111101 : color = 12'he73;
15'b0000101010100111110 : color = 12'he73;
15'b0000101010100111111 : color = 12'he73;
15'b0000101010101000000 : color = 12'he73;
15'b0000101010101000001 : color = 12'he73;
15'b0000101010101000010 : color = 12'he73;
15'b0000101010101000011 : color = 12'he73;
15'b0000101010101000100 : color = 12'he73;
15'b0000101010101000101 : color = 12'he73;
15'b0000101010101000110 : color = 12'he73;
15'b0000101010101000111 : color = 12'he73;
15'b0000101010101001000 : color = 12'he73;
15'b0000101010101001001 : color = 12'he73;
15'b0000101010101001010 : color = 12'he73;
15'b0000101010101001011 : color = 12'he73;
15'b0000101010101001100 : color = 12'he73;
15'b0000101010101001101 : color = 12'he73;
15'b0000101010101001110 : color = 12'he73;
15'b0000101010101001111 : color = 12'he73;
15'b0000101010101010000 : color = 12'he73;
15'b0000101010101010001 : color = 12'he73;
15'b0000101010101010010 : color = 12'he73;
15'b0000101010101010011 : color = 12'he73;
15'b0000101010101010100 : color = 12'he73;
15'b0000101010101010101 : color = 12'he73;
15'b0000101010101010110 : color = 12'he73;
15'b0000101010101010111 : color = 12'he73;
15'b0000101010101011000 : color = 12'he73;
15'b0000101010101011001 : color = 12'he73;
15'b0000101010101011010 : color = 12'he73;
15'b0000101010101011011 : color = 12'he73;
15'b0000101010101011100 : color = 12'he73;
15'b0000101010101011101 : color = 12'he73;
15'b0000101010101011110 : color = 12'he73;
15'b0000101010101011111 : color = 12'he73;
15'b0000101010101100000 : color = 12'he73;
15'b0000101010101100001 : color = 12'he73;
15'b0000101010101100010 : color = 12'he73;
15'b0000101010101100011 : color = 12'he73;
15'b0000101010101100100 : color = 12'he73;
15'b0000101010101100101 : color = 12'he73;
15'b0000101010101100110 : color = 12'he73;
15'b0000101010101100111 : color = 12'he73;
15'b0000101010101101000 : color = 12'he73;
15'b0000101010101101001 : color = 12'he73;
15'b0000101010101101010 : color = 12'he73;
15'b0000101010101101011 : color = 12'he73;
15'b0000101010101101100 : color = 12'he73;
15'b0000101010101101101 : color = 12'he73;
15'b0000101010101101110 : color = 12'he73;
15'b0000101010101101111 : color = 12'he73;
15'b0000101010101110000 : color = 12'he73;
15'b0000101010101110001 : color = 12'he73;
15'b0000101010101110010 : color = 12'he73;
15'b0000101010101110011 : color = 12'he73;
15'b0000101010101110100 : color = 12'he73;
15'b0000101010101110101 : color = 12'he73;
15'b0000101010101110110 : color = 12'he73;
15'b0000101010101110111 : color = 12'he73;
15'b0000101010101111000 : color = 12'he73;
15'b0000101010101111001 : color = 12'he73;
15'b0000101010101111010 : color = 12'he73;
15'b0000101010101111011 : color = 12'he73;
15'b0000101010101111100 : color = 12'he73;
15'b0000101010101111101 : color = 12'he73;
15'b0000101010101111110 : color = 12'he73;
15'b0000101010101111111 : color = 12'he73;
15'b0000101010110000000 : color = 12'he73;
15'b0000101010110000001 : color = 12'he73;
15'b0000101010110000010 : color = 12'he73;
15'b0000101010110000011 : color = 12'he73;
15'b0000101010110000100 : color = 12'he73;
15'b0000101010110000101 : color = 12'he73;
15'b0000101010110000110 : color = 12'he73;
15'b0000101010110000111 : color = 12'he73;
15'b0000101010110001000 : color = 12'he73;
15'b0000101010110001001 : color = 12'he73;
15'b0000101010110001010 : color = 12'he73;
15'b0000101010110001011 : color = 12'he73;
15'b0000101010110001100 : color = 12'he73;
15'b0000101010110001101 : color = 12'he73;
15'b0000101010110001110 : color = 12'he73;
15'b0000101010110001111 : color = 12'he73;
15'b0000101010110010000 : color = 12'he73;
15'b0000101010110010001 : color = 12'he73;
15'b0000101010110010010 : color = 12'he73;
15'b0000101010110010011 : color = 12'he73;
15'b0000101010110010100 : color = 12'he73;
15'b0000101010110010101 : color = 12'he73;
15'b0000101010110010110 : color = 12'he73;
15'b0000101010110010111 : color = 12'he73;
15'b0000101010110011000 : color = 12'he73;
15'b0000101010110011001 : color = 12'he73;
15'b0000101010110011010 : color = 12'he73;
15'b0000101010110011011 : color = 12'he73;
15'b0000101010110011100 : color = 12'he73;
15'b0000101010110011101 : color = 12'he73;
15'b0000101010110011110 : color = 12'he73;
15'b0000101010110011111 : color = 12'he73;
15'b0000101010110100000 : color = 12'he73;
15'b0000101010110100001 : color = 12'he73;
15'b0000101010110100010 : color = 12'he73;
15'b0000101010110100011 : color = 12'he73;
15'b0000101010110100100 : color = 12'he73;
15'b0000101010110100101 : color = 12'he73;
15'b0000101010110100110 : color = 12'he73;
15'b0000101010110100111 : color = 12'he73;
15'b0000101010110101000 : color = 12'he73;
15'b0000101010110101001 : color = 12'he73;
15'b0000101010110101010 : color = 12'he73;
15'b0000101010110101011 : color = 12'he73;
15'b0000101010110101100 : color = 12'he73;
15'b0000101010110101101 : color = 12'he73;
15'b0000101010110101110 : color = 12'he73;
15'b0000101010110101111 : color = 12'he73;
15'b0000101010110110000 : color = 12'he73;
15'b0000101010110110001 : color = 12'he73;
15'b0000101010110110010 : color = 12'he73;
15'b0000101010110110011 : color = 12'he73;
15'b0000101010110110100 : color = 12'he73;
15'b0000101010110110101 : color = 12'he73;
15'b0000101010110110110 : color = 12'he73;
15'b0000101010110110111 : color = 12'he73;
15'b0000101010110111000 : color = 12'he73;
15'b0000101010110111001 : color = 12'he73;
15'b0000101010110111010 : color = 12'he73;
15'b0000101010110111011 : color = 12'he73;
15'b0000101010110111100 : color = 12'he73;
15'b0000101010110111101 : color = 12'he73;
15'b0000101010110111110 : color = 12'he73;
15'b0000101010110111111 : color = 12'he73;
15'b0000101010111000000 : color = 12'he73;
15'b0000101010111000001 : color = 12'he73;
15'b0000101010111000010 : color = 12'he73;
15'b0000101010111000011 : color = 12'he73;
15'b0000101010111000100 : color = 12'he73;
15'b0000101010111000101 : color = 12'he73;
15'b0000101010111000110 : color = 12'he73;
15'b0000101010111000111 : color = 12'he73;
15'b0000101010111001000 : color = 12'he73;
15'b0000101010111001001 : color = 12'he73;
15'b0000101010111001010 : color = 12'he73;
15'b0000101010111001011 : color = 12'he73;
15'b0000101010111001100 : color = 12'he73;
15'b0000101010111001101 : color = 12'he73;
15'b0000101010111001110 : color = 12'he73;
15'b0000101010111001111 : color = 12'he73;
15'b0000101010111010000 : color = 12'he73;
15'b0000101010111010001 : color = 12'he73;
15'b0000101010111010010 : color = 12'he73;
15'b0000101010111010011 : color = 12'he73;
15'b0000101010111010100 : color = 12'he73;
15'b0000101010111010101 : color = 12'he73;
15'b0000101010111010110 : color = 12'he73;
15'b0000101010111010111 : color = 12'he73;
15'b0000101010111011000 : color = 12'he73;
15'b0000101010111011001 : color = 12'he73;
15'b0000101010111011010 : color = 12'he73;
15'b0000101010111011011 : color = 12'he73;
15'b0000101010111011100 : color = 12'he73;
15'b0000101010111011101 : color = 12'he73;
15'b0000101010111011110 : color = 12'he73;
15'b0000101010111011111 : color = 12'he73;
15'b0000101010111100000 : color = 12'he73;
15'b0000101010111100001 : color = 12'he73;
15'b0000101010111100010 : color = 12'he73;
15'b0000101010111100011 : color = 12'he73;
15'b0000101010111100100 : color = 12'he73;
15'b0000101010111100101 : color = 12'he73;
15'b0000101010111100110 : color = 12'he73;
15'b0000101010111100111 : color = 12'he73;
15'b0000101010111101000 : color = 12'he73;
15'b0000101010111101001 : color = 12'he73;
15'b0000101010111101010 : color = 12'he73;
15'b0000101010111101011 : color = 12'he73;
15'b0000101010111101100 : color = 12'he73;
15'b0000101010111101101 : color = 12'he73;
15'b0000101010111101110 : color = 12'he73;
15'b0000101010111101111 : color = 12'he73;
15'b0000101010111110000 : color = 12'he73;
15'b0000101010111110001 : color = 12'he73;
15'b0000101010111110010 : color = 12'he73;
15'b0000101010111110011 : color = 12'he73;
15'b0000101010111110100 : color = 12'he73;
15'b0000101010111110101 : color = 12'he73;
15'b0000101010111110110 : color = 12'he73;
15'b0000101010111110111 : color = 12'he73;
15'b0000101010111111000 : color = 12'he73;
15'b0000101010111111001 : color = 12'he73;
15'b0000101010111111010 : color = 12'he73;
15'b0000101010111111011 : color = 12'he73;
15'b0000101010111111100 : color = 12'he73;
15'b0000101010111111101 : color = 12'he73;
15'b0000101010111111110 : color = 12'he73;
15'b0000101010111111111 : color = 12'he73;
15'b0000101011000000000 : color = 12'he73;
15'b0000101011000000001 : color = 12'he73;
15'b0000101011000000010 : color = 12'he73;
15'b0000101011000000011 : color = 12'he73;
15'b0000101011000000100 : color = 12'he73;
15'b0000101011000000101 : color = 12'he73;
15'b0000101011000000110 : color = 12'he73;
15'b0000101011000000111 : color = 12'he73;
15'b0000101011000001000 : color = 12'he73;
15'b0000101011000001001 : color = 12'he73;
15'b0000101011000001010 : color = 12'he73;
15'b0000101011000001011 : color = 12'he73;
15'b0000101011000001100 : color = 12'he73;
15'b0000101011000001101 : color = 12'he73;
15'b0000101011000001110 : color = 12'he73;
15'b0000101011000001111 : color = 12'he73;
15'b0000101011000010000 : color = 12'he73;
15'b0000101011000010001 : color = 12'he73;
15'b0000101011000010010 : color = 12'he73;
15'b0000101011000010011 : color = 12'he73;
15'b0000101011000010100 : color = 12'he73;
15'b0000101011000010101 : color = 12'he73;
15'b0000101011000010110 : color = 12'he73;
15'b0000101011000010111 : color = 12'he73;
15'b0000101011000011000 : color = 12'he73;
15'b0000101011000011001 : color = 12'he73;
15'b0000101011000011010 : color = 12'he73;
15'b0000101011000011011 : color = 12'he73;
15'b0000101011000011100 : color = 12'he73;
15'b0000101011000011101 : color = 12'he73;
15'b0000101011000011110 : color = 12'he73;
15'b0000101011000011111 : color = 12'he73;
15'b0000101011000100000 : color = 12'he73;
15'b0000101011000100001 : color = 12'he73;
15'b0000101011000100010 : color = 12'he73;
15'b0000101011000100011 : color = 12'he73;
15'b0000101011000100100 : color = 12'he73;
15'b0000101011000100101 : color = 12'he73;
15'b0000101011000100110 : color = 12'he73;
15'b0000101011000100111 : color = 12'he73;
15'b0000101011000101000 : color = 12'he73;
15'b0000101011000101001 : color = 12'he73;
15'b0000101011000101010 : color = 12'he73;
15'b0000101011000101011 : color = 12'he73;
15'b0000101011000101100 : color = 12'he73;
15'b0000101011000101101 : color = 12'he73;
15'b0000101011000101110 : color = 12'he73;
15'b0000101011000101111 : color = 12'he73;
15'b0000101011000110000 : color = 12'he73;
15'b0000101011000110001 : color = 12'he73;
15'b0000101011000110010 : color = 12'he73;
15'b0000101011000110011 : color = 12'he73;
15'b0000101011000110100 : color = 12'he73;
15'b0000101011000110101 : color = 12'he73;
15'b0000101011000110110 : color = 12'he73;
15'b0000101011000110111 : color = 12'he73;
15'b0000101011000111000 : color = 12'he73;
15'b0000101011000111001 : color = 12'he73;
15'b0000101011000111010 : color = 12'he73;
15'b0000101011000111011 : color = 12'he73;
15'b0000101011000111100 : color = 12'he73;
15'b0000101011000111101 : color = 12'he73;
15'b0000101011000111110 : color = 12'he73;
15'b0000101011000111111 : color = 12'he73;
15'b0000101011001000000 : color = 12'he73;
15'b0000101011001000001 : color = 12'he73;
15'b0000101011001000010 : color = 12'he73;
15'b0000101011001000011 : color = 12'he73;
15'b0000101011001000100 : color = 12'he73;
15'b0000101011001000101 : color = 12'he73;
15'b0000101011001000110 : color = 12'he73;
15'b0000101011001000111 : color = 12'he73;
15'b0000101011001001000 : color = 12'he73;
15'b0000101011001001001 : color = 12'he73;
15'b0000101011001001010 : color = 12'he73;
15'b0000101011001001011 : color = 12'he73;
15'b0000101011001001100 : color = 12'he73;
15'b0000101011001001101 : color = 12'he73;
15'b0000101011001001110 : color = 12'he73;
15'b0000101011001001111 : color = 12'he73;
15'b0000101011001010000 : color = 12'he73;
15'b0000101011001010001 : color = 12'he73;
15'b0000101010010010000 : color = 12'he73;
15'b0000101010010010001 : color = 12'he73;
15'b0000101010010010010 : color = 12'he73;
15'b0000101010010010011 : color = 12'he73;
15'b0000101010010010100 : color = 12'he73;
15'b0000101010010010101 : color = 12'he73;
15'b0000101010010010110 : color = 12'he73;
15'b0000101010010010111 : color = 12'he73;
15'b0000101010010011000 : color = 12'he73;
15'b0000101010010011001 : color = 12'he73;
15'b0000101010010011010 : color = 12'he73;
15'b0000101010010011011 : color = 12'he73;
15'b0000101010010011100 : color = 12'he73;
15'b0000101010010011101 : color = 12'he73;
15'b0000101010010011110 : color = 12'he73;
15'b0000101010010011111 : color = 12'he73;
15'b0000101010010100000 : color = 12'he73;
15'b0000101010010100001 : color = 12'he73;
15'b0000101010010100010 : color = 12'he73;
15'b0000101010010100011 : color = 12'he73;
15'b0000101010010100100 : color = 12'he73;
15'b0000101010010100101 : color = 12'he73;
15'b0000101010010100110 : color = 12'he73;
15'b0000101010010100111 : color = 12'he73;
15'b0000101010010101000 : color = 12'he73;
15'b0000101010010101001 : color = 12'he73;
15'b0000101010010101010 : color = 12'he73;
15'b0000101010010101011 : color = 12'he73;
15'b0000101010010101100 : color = 12'he73;
15'b0000101010010101101 : color = 12'he73;
15'b0000101010010101110 : color = 12'he73;
15'b0000101010010101111 : color = 12'he73;
15'b0000101010010110000 : color = 12'he73;
15'b0000101010010110001 : color = 12'he73;
15'b0000101010010110010 : color = 12'he73;
15'b0000101010010110011 : color = 12'he73;
15'b0000101010010110100 : color = 12'he73;
15'b0000101010010110101 : color = 12'he73;
15'b0000101010010110110 : color = 12'he73;
15'b0000101010010110111 : color = 12'he73;
15'b0000101010010111000 : color = 12'he73;
15'b0000101010010111001 : color = 12'he73;
15'b0000101010010111010 : color = 12'he73;
15'b0000101010010111011 : color = 12'he73;
15'b0000101010010111100 : color = 12'he73;
15'b0000101010010111101 : color = 12'he73;
15'b0000101010010111110 : color = 12'he73;
15'b0000101010010111111 : color = 12'he73;
15'b0000101010011000000 : color = 12'he73;
15'b0000101010011000001 : color = 12'he73;
15'b0000101010011000010 : color = 12'he73;
15'b0000101010011000011 : color = 12'he73;
15'b0000101010011000100 : color = 12'he73;
15'b0000101010011000101 : color = 12'he73;
15'b0000101010011000110 : color = 12'he73;
15'b0000101010011000111 : color = 12'he73;
15'b0000101010011001000 : color = 12'he73;
15'b0000101010011001001 : color = 12'he73;
15'b0000101010011001010 : color = 12'he73;
15'b0000101010011001011 : color = 12'he73;
15'b0000101010011001100 : color = 12'he73;
15'b0000101010011001101 : color = 12'he73;
15'b0000101010011001110 : color = 12'he73;
15'b0000101010011001111 : color = 12'he73;
15'b0000101010011010000 : color = 12'he73;
15'b0000101010011010001 : color = 12'he73;
15'b0000101010011010010 : color = 12'he73;
15'b0000101010011010011 : color = 12'he73;
15'b0000101010011010100 : color = 12'he73;
15'b0000101010011010101 : color = 12'he73;
15'b0000101010011010110 : color = 12'he73;
15'b0000101010011010111 : color = 12'he73;
15'b0000101010011011000 : color = 12'he73;
15'b0000101010011011001 : color = 12'he73;
15'b0000101010011011010 : color = 12'he73;
15'b0000101010011011011 : color = 12'he73;
15'b0000101010011011100 : color = 12'he73;
15'b0000101010011011101 : color = 12'he73;
15'b0000101010011011110 : color = 12'he73;
15'b0000101010011011111 : color = 12'he73;
15'b0000101010011100000 : color = 12'he73;
15'b0000101010011100001 : color = 12'he73;
15'b0000101010011100010 : color = 12'he73;
15'b0000101010011100011 : color = 12'he73;
15'b0000101010011100100 : color = 12'he73;
15'b0000101010011100101 : color = 12'he73;
15'b0000101010011100110 : color = 12'he73;
15'b0000101010011100111 : color = 12'he73;
15'b0000101010011101000 : color = 12'he73;
15'b0000101010011101001 : color = 12'he73;
15'b0000101010011101010 : color = 12'he73;
15'b0000101010011101011 : color = 12'he73;
15'b0000101010011101100 : color = 12'he73;
15'b0000101010011101101 : color = 12'he73;
15'b0000101010011101110 : color = 12'he73;
15'b0000101010011101111 : color = 12'he73;
15'b0000101010011110000 : color = 12'he73;
15'b0000101010011110001 : color = 12'he73;
15'b0000101010011110010 : color = 12'he73;
15'b0000101010011110011 : color = 12'he73;
15'b0000101010011110100 : color = 12'he73;
15'b0000101010011110101 : color = 12'he73;
15'b0000101010011110110 : color = 12'he73;
15'b0000101010011110111 : color = 12'he73;
15'b0000101010011111000 : color = 12'he73;
15'b0000101010011111001 : color = 12'he73;
15'b0000101010011111010 : color = 12'he73;
15'b0000101010011111011 : color = 12'he73;
15'b0000101010011111100 : color = 12'he73;
15'b0000101010011111101 : color = 12'he73;
15'b0000101010011111110 : color = 12'he73;
15'b0000101010011111111 : color = 12'he73;
15'b0000101010100000000 : color = 12'he73;
15'b0000101010100000001 : color = 12'he73;
15'b0000101010100000010 : color = 12'he73;
15'b0000101010100000011 : color = 12'he73;
15'b0000101010100000100 : color = 12'he73;
15'b0000101010100000101 : color = 12'he73;
15'b0000101010100000110 : color = 12'he73;
15'b0000101010100000111 : color = 12'he73;
15'b0000101010100001000 : color = 12'he73;
15'b0000101010100001001 : color = 12'he73;
15'b0000101010100001010 : color = 12'he73;
15'b0000101010100001011 : color = 12'he73;
15'b0000101010100001100 : color = 12'he73;
15'b0000101010100001101 : color = 12'he73;
15'b0000101010100001110 : color = 12'he73;
15'b0000101010100001111 : color = 12'he73;
15'b0000101010100010000 : color = 12'he73;
15'b0000101010100010001 : color = 12'he73;
15'b0000101010100010010 : color = 12'he73;
15'b0000101010100010011 : color = 12'he73;
15'b0000101010100010100 : color = 12'he73;
15'b0000101010100010101 : color = 12'he73;
15'b0000101010100010110 : color = 12'he73;
15'b0000101010100010111 : color = 12'he73;
15'b0000101010100011000 : color = 12'he73;
15'b0000101010100011001 : color = 12'he73;
15'b0000101010100011010 : color = 12'he73;
15'b0000101010100011011 : color = 12'he73;
15'b0000101010100011100 : color = 12'he73;
15'b0000101010100011101 : color = 12'he73;
15'b0000101010100011110 : color = 12'he73;
15'b0000101010100011111 : color = 12'he73;
15'b0000101010100100000 : color = 12'he73;
15'b0000101010100100001 : color = 12'he73;
15'b0000101010100100010 : color = 12'he73;
15'b0000101010100100011 : color = 12'he73;
15'b0000101010100100100 : color = 12'he73;
15'b0000101010100100101 : color = 12'he73;
15'b0000101010100100110 : color = 12'he73;
15'b0000101010100100111 : color = 12'he73;
15'b0000101010100101000 : color = 12'he73;
15'b0000101010100101001 : color = 12'he73;
15'b0000101010100101010 : color = 12'he73;
15'b0000101010100101011 : color = 12'he73;
15'b0000101010100101100 : color = 12'he73;
15'b0000101010100101101 : color = 12'he73;
15'b0000101010100101110 : color = 12'he73;
15'b0000101010100101111 : color = 12'he73;
15'b0000101010100110000 : color = 12'he73;
15'b0000101010100110001 : color = 12'he73;
15'b0000101010100110010 : color = 12'he73;
15'b0000101010100110011 : color = 12'he73;
15'b0000101010100110100 : color = 12'he73;
15'b0000101010100110101 : color = 12'he73;
15'b0000101010100110110 : color = 12'he73;
15'b0000101010100110111 : color = 12'he73;
15'b0000101010100111000 : color = 12'he73;
15'b0000101010100111001 : color = 12'he73;
15'b0000101010100111010 : color = 12'he73;
15'b0000101010100111011 : color = 12'he73;
15'b0000101010100111100 : color = 12'he73;
15'b0000101010100111101 : color = 12'he73;
15'b0000101010100111110 : color = 12'he73;
15'b0000101010100111111 : color = 12'he73;
15'b0000101010101000000 : color = 12'he73;
15'b0000101010101000001 : color = 12'he73;
15'b0000101010101000010 : color = 12'he73;
15'b0000101010101000011 : color = 12'he73;
15'b0000101010101000100 : color = 12'he73;
15'b0000101010101000101 : color = 12'he73;
15'b0000101010101000110 : color = 12'he73;
15'b0000101010101000111 : color = 12'he73;
15'b0000101010101001000 : color = 12'he73;
15'b0000101010101001001 : color = 12'he73;
15'b0000101010101001010 : color = 12'he73;
15'b0000101010101001011 : color = 12'he73;
15'b0000101010101001100 : color = 12'he73;
15'b0000101010101001101 : color = 12'he73;
15'b0000101010101001110 : color = 12'he73;
15'b0000101010101001111 : color = 12'he73;
15'b0000101010101010000 : color = 12'he73;
15'b0000101010101010001 : color = 12'he73;
15'b0000101010101010010 : color = 12'he73;
15'b0000101010101010011 : color = 12'he73;
15'b0000101010101010100 : color = 12'he73;
15'b0000101010101010101 : color = 12'he73;
15'b0000101010101010110 : color = 12'he73;
15'b0000101010101010111 : color = 12'he73;
15'b0000101010101011000 : color = 12'he73;
15'b0000101010101011001 : color = 12'he73;
15'b0000101010101011010 : color = 12'he73;
15'b0000101010101011011 : color = 12'he73;
15'b0000101010101011100 : color = 12'he73;
15'b0000101010101011101 : color = 12'he73;
15'b0000101010101011110 : color = 12'he73;
15'b0000101010101011111 : color = 12'he73;
15'b0000101010101100000 : color = 12'he73;
15'b0000101010101100001 : color = 12'he73;
15'b0000101010101100010 : color = 12'he73;
15'b0000101010101100011 : color = 12'he73;
15'b0000101010101100100 : color = 12'he73;
15'b0000101010101100101 : color = 12'he73;
15'b0000101010101100110 : color = 12'he73;
15'b0000101010101100111 : color = 12'he73;
15'b0000101010101101000 : color = 12'he73;
15'b0000101010101101001 : color = 12'he73;
15'b0000101010101101010 : color = 12'he73;
15'b0000101010101101011 : color = 12'he73;
15'b0000101010101101100 : color = 12'he73;
15'b0000101010101101101 : color = 12'he73;
15'b0000101010101101110 : color = 12'he73;
15'b0000101010101101111 : color = 12'he73;
15'b0000101010101110000 : color = 12'he73;
15'b0000101010101110001 : color = 12'he73;
15'b0000101010101110010 : color = 12'he73;
15'b0000101010101110011 : color = 12'he73;
15'b0000101010101110100 : color = 12'he73;
15'b0000101010101110101 : color = 12'he73;
15'b0000101010101110110 : color = 12'he73;
15'b0000101010101110111 : color = 12'he73;
15'b0000101010101111000 : color = 12'he73;
15'b0000101010101111001 : color = 12'he73;
15'b0000101010101111010 : color = 12'he73;
15'b0000101010101111011 : color = 12'he73;
15'b0000101010101111100 : color = 12'he73;
15'b0000101010101111101 : color = 12'he73;
15'b0000101010101111110 : color = 12'he73;
15'b0000101010101111111 : color = 12'he73;
15'b0000101010110000000 : color = 12'he73;
15'b0000101010110000001 : color = 12'he73;
15'b0000101010110000010 : color = 12'he73;
15'b0000101010110000011 : color = 12'he73;
15'b0000101010110000100 : color = 12'he73;
15'b0000101010110000101 : color = 12'he73;
15'b0000101010110000110 : color = 12'he73;
15'b0000101010110000111 : color = 12'he73;
15'b0000101010110001000 : color = 12'he73;
15'b0000101010110001001 : color = 12'he73;
15'b0000101010110001010 : color = 12'he73;
15'b0000101010110001011 : color = 12'he73;
15'b0000101010110001100 : color = 12'he73;
15'b0000101010110001101 : color = 12'he73;
15'b0000101010110001110 : color = 12'he73;
15'b0000101010110001111 : color = 12'he73;
15'b0000101010110010000 : color = 12'he73;
15'b0000101010110010001 : color = 12'he73;
15'b0000101010110010010 : color = 12'he73;
15'b0000101010110010011 : color = 12'he73;
15'b0000101010110010100 : color = 12'he73;
15'b0000101010110010101 : color = 12'he73;
15'b0000101010110010110 : color = 12'he73;
15'b0000101010110010111 : color = 12'he73;
15'b0000101010110011000 : color = 12'he73;
15'b0000101010110011001 : color = 12'he73;
15'b0000101010110011010 : color = 12'he73;
15'b0000101010110011011 : color = 12'he73;
15'b0000101010110011100 : color = 12'he73;
15'b0000101010110011101 : color = 12'he73;
15'b0000101010110011110 : color = 12'he73;
15'b0000101010110011111 : color = 12'he73;
15'b0000101010110100000 : color = 12'he73;
15'b0000101010110100001 : color = 12'he73;
15'b0000101010110100010 : color = 12'he73;
15'b0000101010110100011 : color = 12'he73;
15'b0000101010110100100 : color = 12'he73;
15'b0000101010110100101 : color = 12'he73;
15'b0000101010110100110 : color = 12'he73;
15'b0000101010110100111 : color = 12'he73;
15'b0000101010110101000 : color = 12'he73;
15'b0000101010110101001 : color = 12'he73;
15'b0000101010110101010 : color = 12'he73;
15'b0000101010110101011 : color = 12'he73;
15'b0000101010110101100 : color = 12'he73;
15'b0000101010110101101 : color = 12'he73;
15'b0000101010110101110 : color = 12'he73;
15'b0000101010110101111 : color = 12'he73;
15'b0000101010110110000 : color = 12'he73;
15'b0000101010110110001 : color = 12'he73;
15'b0000101010110110010 : color = 12'he73;
15'b0000101010110110011 : color = 12'he73;
15'b0000101010110110100 : color = 12'he73;
15'b0000101010110110101 : color = 12'he73;
15'b0000101010110110110 : color = 12'he73;
15'b0000101010110110111 : color = 12'he73;
15'b0000101010110111000 : color = 12'he73;
15'b0000101010110111001 : color = 12'he73;
15'b0000101010110111010 : color = 12'he73;
15'b0000101010110111011 : color = 12'he73;
15'b0000101010110111100 : color = 12'he73;
15'b0000101010110111101 : color = 12'he73;
15'b0000101010110111110 : color = 12'he73;
15'b0000101010110111111 : color = 12'he73;
15'b0000101010111000000 : color = 12'he73;
15'b0000101010111000001 : color = 12'he73;
15'b0000101010111000010 : color = 12'he73;
15'b0000101010111000011 : color = 12'he73;
15'b0000101010111000100 : color = 12'he73;
15'b0000101010111000101 : color = 12'he73;
15'b0000101010111000110 : color = 12'he73;
15'b0000101010111000111 : color = 12'he73;
15'b0000101010111001000 : color = 12'he73;
15'b0000101010111001001 : color = 12'he73;
15'b0000101010111001010 : color = 12'he73;
15'b0000101010111001011 : color = 12'he73;
15'b0000101010111001100 : color = 12'he73;
15'b0000101010111001101 : color = 12'he73;
15'b0000101010111001110 : color = 12'he73;
15'b0000101010111001111 : color = 12'he73;
15'b0000101010111010000 : color = 12'he73;
15'b0000101010111010001 : color = 12'he73;
15'b0000101010111010010 : color = 12'he73;
15'b0000101010111010011 : color = 12'he73;
15'b0000101010111010100 : color = 12'he73;
15'b0000101010111010101 : color = 12'he73;
15'b0000101010111010110 : color = 12'he73;
15'b0000101010111010111 : color = 12'he73;
15'b0000101010111011000 : color = 12'he73;
15'b0000101010111011001 : color = 12'he73;
15'b0000101010111011010 : color = 12'he73;
15'b0000101010111011011 : color = 12'he73;
15'b0000101010111011100 : color = 12'he73;
15'b0000101010111011101 : color = 12'he73;
15'b0000101010111011110 : color = 12'he73;
15'b0000101010111011111 : color = 12'he73;
15'b0000101010111100000 : color = 12'he73;
15'b0000101010111100001 : color = 12'he73;
15'b0000101010111100010 : color = 12'he73;
15'b0000101010111100011 : color = 12'he73;
15'b0000101010111100100 : color = 12'he73;
15'b0000101010111100101 : color = 12'he73;
15'b0000101010111100110 : color = 12'he73;
15'b0000101010111100111 : color = 12'he73;
15'b0000101010111101000 : color = 12'he73;
15'b0000101010111101001 : color = 12'he73;
15'b0000101010111101010 : color = 12'he73;
15'b0000101010111101011 : color = 12'he73;
15'b0000101010111101100 : color = 12'he73;
15'b0000101010111101101 : color = 12'he73;
15'b0000101010111101110 : color = 12'he73;
15'b0000101010111101111 : color = 12'he73;
15'b0000101010111110000 : color = 12'he73;
15'b0000101010111110001 : color = 12'he73;
15'b0000101010111110010 : color = 12'he73;
15'b0000101010111110011 : color = 12'he73;
15'b0000101010111110100 : color = 12'he73;
15'b0000101010111110101 : color = 12'he73;
15'b0000101010111110110 : color = 12'he73;
15'b0000101010111110111 : color = 12'he73;
15'b0000101010111111000 : color = 12'he73;
15'b0000101010111111001 : color = 12'he73;
15'b0000101010111111010 : color = 12'he73;
15'b0000101010111111011 : color = 12'he73;
15'b0000101010111111100 : color = 12'he73;
15'b0000101010111111101 : color = 12'he73;
15'b0000101010111111110 : color = 12'he73;
15'b0000101010111111111 : color = 12'he73;
15'b0000101011000000000 : color = 12'he73;
15'b0000101011000000001 : color = 12'he73;
15'b0000101011000000010 : color = 12'he73;
15'b0000101011000000011 : color = 12'he73;
15'b0000101011000000100 : color = 12'he73;
15'b0000101011000000101 : color = 12'he73;
15'b0000101011000000110 : color = 12'he73;
15'b0000101011000000111 : color = 12'he73;
15'b0000101011000001000 : color = 12'he73;
15'b0000101011000001001 : color = 12'he73;
15'b0000101011000001010 : color = 12'he73;
15'b0000101011000001011 : color = 12'he73;
15'b0000101011000001100 : color = 12'he73;
15'b0000101011000001101 : color = 12'he73;
15'b0000101011000001110 : color = 12'he73;
15'b0000101011000001111 : color = 12'he73;
15'b0000101011000010000 : color = 12'he73;
15'b0000101011000010001 : color = 12'he73;
15'b0000101011000010010 : color = 12'he73;
15'b0000101011000010011 : color = 12'he73;
15'b0000101011000010100 : color = 12'he73;
15'b0000101011000010101 : color = 12'he73;
15'b0000101011000010110 : color = 12'he73;
15'b0000101011000010111 : color = 12'he73;
15'b0000101011000011000 : color = 12'he73;
15'b0000101011000011001 : color = 12'he73;
15'b0000101011000011010 : color = 12'he73;
15'b0000101011000011011 : color = 12'he73;
15'b0000101011000011100 : color = 12'he73;
15'b0000101011000011101 : color = 12'he73;
15'b0000101011000011110 : color = 12'he73;
15'b0000101011000011111 : color = 12'he73;
15'b0000101011000100000 : color = 12'he73;
15'b0000101011000100001 : color = 12'he73;
15'b0000101011000100010 : color = 12'he73;
15'b0000101011000100011 : color = 12'he73;
15'b0000101011000100100 : color = 12'he73;
15'b0000101011000100101 : color = 12'he73;
15'b0000101011000100110 : color = 12'he73;
15'b0000101011000100111 : color = 12'he73;
15'b0000101011000101000 : color = 12'he73;
15'b0000101011000101001 : color = 12'he73;
15'b0000101011000101010 : color = 12'he73;
15'b0000101011000101011 : color = 12'he73;
15'b0000101011000101100 : color = 12'he73;
15'b0000101011000101101 : color = 12'he73;
15'b0000101011000101110 : color = 12'he73;
15'b0000101011000101111 : color = 12'he73;
15'b0000101011000110000 : color = 12'he73;
15'b0000101011000110001 : color = 12'he73;
15'b0000101011000110010 : color = 12'he73;
15'b0000101011000110011 : color = 12'he73;
15'b0000101011000110100 : color = 12'he73;
15'b0000101011000110101 : color = 12'he73;
15'b0000101011000110110 : color = 12'he73;
15'b0000101011000110111 : color = 12'he73;
15'b0000101011000111000 : color = 12'he73;
15'b0000101011000111001 : color = 12'he73;
15'b0000101011000111010 : color = 12'he73;
15'b0000101011000111011 : color = 12'he73;
15'b0000101011000111100 : color = 12'he73;
15'b0000101011000111101 : color = 12'he73;
15'b0000101011000111110 : color = 12'he73;
15'b0000101011000111111 : color = 12'he73;
15'b0000101011001000000 : color = 12'he73;
15'b0000101011001000001 : color = 12'he73;
15'b0000101011001000010 : color = 12'he73;
15'b0000101011001000011 : color = 12'he73;
15'b0000101011001000100 : color = 12'he73;
15'b0000101011001000101 : color = 12'he73;
15'b0000101011001000110 : color = 12'he73;
15'b0000101011001000111 : color = 12'he73;
15'b0000101011001001000 : color = 12'he73;
15'b0000101011001001001 : color = 12'he73;
15'b0000101011001001010 : color = 12'he73;
15'b0000101011001001011 : color = 12'he73;
15'b0000101011001001100 : color = 12'he73;
15'b0000101011001001101 : color = 12'he73;
15'b0000101011001001110 : color = 12'he73;
15'b0000101011001001111 : color = 12'he73;
15'b0000101011001010000 : color = 12'he73;
15'b0000101011001010001 : color = 12'he73;
15'b0000101011001010010 : color = 12'he73;
15'b0000101011001010011 : color = 12'he73;
15'b0000101011001010100 : color = 12'he73;
15'b0000101011001010101 : color = 12'he73;
15'b0000101011001010110 : color = 12'he73;
15'b0000101011001010111 : color = 12'he73;
15'b0000101011001011000 : color = 12'he73;
15'b0000101011001011001 : color = 12'he73;
15'b0000101011001011010 : color = 12'he73;
15'b0000101011001011011 : color = 12'he73;
15'b0000101011001011100 : color = 12'he73;
15'b0000101011001011101 : color = 12'he73;
15'b0000101011001011110 : color = 12'he73;
15'b0000101011001011111 : color = 12'he73;
15'b0000101011001100000 : color = 12'he73;
15'b0000101011001100001 : color = 12'he73;
15'b0000101011001100010 : color = 12'he73;
15'b0000101011001100011 : color = 12'he73;
15'b0000101011001100100 : color = 12'he73;
15'b0000101011001100101 : color = 12'he73;
15'b0000101011001100110 : color = 12'he73;
15'b0000101011001100111 : color = 12'he73;
15'b0000101011001101000 : color = 12'he73;
15'b0000101011001101001 : color = 12'he73;
15'b0000101011001101010 : color = 12'he73;
15'b0000101011001101011 : color = 12'he73;
15'b0000101011001101100 : color = 12'he73;
15'b0000101011001101101 : color = 12'he73;
15'b0000101011001101110 : color = 12'he73;
15'b0000101011001101111 : color = 12'he73;
15'b0000101011001110000 : color = 12'he73;
15'b0000101011001110001 : color = 12'he73;
15'b0000101011001110010 : color = 12'he73;
15'b0000101011001110011 : color = 12'he73;
15'b0000101011001110100 : color = 12'he73;
15'b0000101011001110101 : color = 12'he73;
15'b0000101011001110110 : color = 12'he73;
15'b0000101011001110111 : color = 12'he73;
15'b0000101011001111000 : color = 12'he73;
15'b0000101011001111001 : color = 12'he73;
15'b0000101011001111010 : color = 12'he73;
15'b0000101010010111001 : color = 12'he73;
15'b0000101010010111010 : color = 12'he73;
15'b0000101010010111011 : color = 12'he73;
15'b0000101010010111100 : color = 12'he73;
15'b0000101010010111101 : color = 12'he73;
15'b0000101010010111110 : color = 12'he73;
15'b0000101010010111111 : color = 12'he73;
15'b0000101010011000000 : color = 12'he73;
15'b0000101010011000001 : color = 12'he73;
15'b0000101010011000010 : color = 12'he73;
15'b0000101010011000011 : color = 12'he73;
15'b0000101010011000100 : color = 12'he73;
15'b0000101010011000101 : color = 12'he73;
15'b0000101010011000110 : color = 12'he73;
15'b0000101010011000111 : color = 12'he73;
15'b0000101010011001000 : color = 12'he73;
15'b0000101010011001001 : color = 12'he73;
15'b0000101010011001010 : color = 12'he73;
15'b0000101010011001011 : color = 12'he73;
15'b0000101010011001100 : color = 12'he73;
15'b0000101010011001101 : color = 12'he73;
15'b0000101010011001110 : color = 12'he73;
15'b0000101010011001111 : color = 12'he73;
15'b0000101010011010000 : color = 12'he73;
15'b0000101010011010001 : color = 12'he73;
15'b0000101010011010010 : color = 12'he73;
15'b0000101010011010011 : color = 12'he73;
15'b0000101010011010100 : color = 12'he73;
15'b0000101010011010101 : color = 12'he73;
15'b0000101010011010110 : color = 12'he73;
15'b0000101010011010111 : color = 12'he73;
15'b0000101010011011000 : color = 12'he73;
15'b0000101010011011001 : color = 12'he73;
15'b0000101010011011010 : color = 12'he73;
15'b0000101010011011011 : color = 12'he73;
15'b0000101010011011100 : color = 12'he73;
15'b0000101010011011101 : color = 12'he73;
15'b0000101010011011110 : color = 12'he73;
15'b0000101010011011111 : color = 12'he73;
15'b0000101010011100000 : color = 12'he73;
15'b0000101010011100001 : color = 12'he73;
15'b0000101010011100010 : color = 12'he73;
15'b0000101010011100011 : color = 12'he73;
15'b0000101010011100100 : color = 12'he73;
15'b0000101010011100101 : color = 12'he73;
15'b0000101010011100110 : color = 12'he73;
15'b0000101010011100111 : color = 12'he73;
15'b0000101010011101000 : color = 12'he73;
15'b0000101010011101001 : color = 12'he73;
15'b0000101010011101010 : color = 12'he73;
15'b0000101010011101011 : color = 12'he73;
15'b0000101010011101100 : color = 12'he73;
15'b0000101010011101101 : color = 12'he73;
15'b0000101010011101110 : color = 12'he73;
15'b0000101010011101111 : color = 12'he73;
15'b0000101010011110000 : color = 12'he73;
15'b0000101010011110001 : color = 12'he73;
15'b0000101010011110010 : color = 12'he73;
15'b0000101010011110011 : color = 12'he73;
15'b0000101010011110100 : color = 12'he73;
15'b0000101010011110101 : color = 12'he73;
15'b0000101010011110110 : color = 12'he73;
15'b0000101010011110111 : color = 12'he73;
15'b0000101010011111000 : color = 12'he73;
15'b0000101010011111001 : color = 12'he73;
15'b0000101010011111010 : color = 12'he73;
15'b0000101010011111011 : color = 12'he73;
15'b0000101010011111100 : color = 12'he73;
15'b0000101010011111101 : color = 12'he73;
15'b0000101010011111110 : color = 12'he73;
15'b0000101010011111111 : color = 12'he73;
15'b0000101010100000000 : color = 12'he73;
15'b0000101010100000001 : color = 12'he73;
15'b0000101010100000010 : color = 12'he73;
15'b0000101010100000011 : color = 12'he73;
15'b0000101010100000100 : color = 12'he73;
15'b0000101010100000101 : color = 12'he73;
15'b0000101010100000110 : color = 12'he73;
15'b0000101010100000111 : color = 12'he73;
15'b0000101010100001000 : color = 12'he73;
15'b0000101010100001001 : color = 12'he73;
15'b0000101010100001010 : color = 12'he73;
15'b0000101010100001011 : color = 12'he73;
15'b0000101010100001100 : color = 12'he73;
15'b0000101010100001101 : color = 12'he73;
15'b0000101010100001110 : color = 12'he73;
15'b0000101010100001111 : color = 12'he73;
15'b0000101010100010000 : color = 12'he73;
15'b0000101010100010001 : color = 12'he73;
15'b0000101010100010010 : color = 12'he73;
15'b0000101010100010011 : color = 12'he73;
15'b0000101010100010100 : color = 12'he73;
15'b0000101010100010101 : color = 12'he73;
15'b0000101010100010110 : color = 12'he73;
15'b0000101010100010111 : color = 12'he73;
15'b0000101010100011000 : color = 12'he73;
15'b0000101010100011001 : color = 12'he73;
15'b0000101010100011010 : color = 12'he73;
15'b0000101010100011011 : color = 12'he73;
15'b0000101010100011100 : color = 12'he73;
15'b0000101010100011101 : color = 12'he73;
15'b0000101010100011110 : color = 12'he73;
15'b0000101010100011111 : color = 12'he73;
15'b0000101010100100000 : color = 12'he73;
15'b0000101010100100001 : color = 12'he73;
15'b0000101010100100010 : color = 12'he73;
15'b0000101010100100011 : color = 12'he73;
15'b0000101010100100100 : color = 12'he73;
15'b0000101010100100101 : color = 12'he73;
15'b0000101010100100110 : color = 12'he73;
15'b0000101010100100111 : color = 12'he73;
15'b0000101010100101000 : color = 12'he73;
15'b0000101010100101001 : color = 12'he73;
15'b0000101010100101010 : color = 12'he73;
15'b0000101010100101011 : color = 12'he73;
15'b0000101010100101100 : color = 12'he73;
15'b0000101010100101101 : color = 12'he73;
15'b0000101010100101110 : color = 12'he73;
15'b0000101010100101111 : color = 12'he73;
15'b0000101010100110000 : color = 12'he73;
15'b0000101010100110001 : color = 12'he73;
15'b0000101010100110010 : color = 12'he73;
15'b0000101010100110011 : color = 12'he73;
15'b0000101010100110100 : color = 12'he73;
15'b0000101010100110101 : color = 12'he73;
15'b0000101010100110110 : color = 12'he73;
15'b0000101010100110111 : color = 12'he73;
15'b0000101010100111000 : color = 12'he73;
15'b0000101010100111001 : color = 12'he73;
15'b0000101010100111010 : color = 12'he73;
15'b0000101010100111011 : color = 12'he73;
15'b0000101010100111100 : color = 12'he73;
15'b0000101010100111101 : color = 12'he73;
15'b0000101010100111110 : color = 12'he73;
15'b0000101010100111111 : color = 12'he73;
15'b0000101010101000000 : color = 12'he73;
15'b0000101010101000001 : color = 12'he73;
15'b0000101010101000010 : color = 12'he73;
15'b0000101010101000011 : color = 12'he73;
15'b0000101010101000100 : color = 12'he73;
15'b0000101010101000101 : color = 12'he73;
15'b0000101010101000110 : color = 12'he73;
15'b0000101010101000111 : color = 12'he73;
15'b0000101010101001000 : color = 12'he73;
15'b0000101010101001001 : color = 12'he73;
15'b0000101010101001010 : color = 12'he73;
15'b0000101010101001011 : color = 12'he73;
15'b0000101010101001100 : color = 12'he73;
15'b0000101010101001101 : color = 12'he73;
15'b0000101010101001110 : color = 12'he73;
15'b0000101010101001111 : color = 12'he73;
15'b0000101010101010000 : color = 12'he73;
15'b0000101010101010001 : color = 12'he73;
15'b0000101010101010010 : color = 12'he73;
15'b0000101010101010011 : color = 12'he73;
15'b0000101010101010100 : color = 12'he73;
15'b0000101010101010101 : color = 12'he73;
15'b0000101010101010110 : color = 12'he73;
15'b0000101010101010111 : color = 12'he73;
15'b0000101010101011000 : color = 12'he73;
15'b0000101010101011001 : color = 12'he73;
15'b0000101010101011010 : color = 12'he73;
15'b0000101010101011011 : color = 12'he73;
15'b0000101010101011100 : color = 12'he73;
15'b0000101010101011101 : color = 12'he73;
15'b0000101010101011110 : color = 12'he73;
15'b0000101010101011111 : color = 12'he73;
15'b0000101010101100000 : color = 12'he73;
15'b0000101010101100001 : color = 12'he73;
15'b0000101010101100010 : color = 12'he73;
15'b0000101010101100011 : color = 12'he73;
15'b0000101010101100100 : color = 12'he73;
15'b0000101010101100101 : color = 12'he73;
15'b0000101010101100110 : color = 12'he73;
15'b0000101010101100111 : color = 12'he73;
15'b0000101010101101000 : color = 12'he73;
15'b0000101010101101001 : color = 12'he73;
15'b0000101010101101010 : color = 12'he73;
15'b0000101010101101011 : color = 12'he73;
15'b0000101010101101100 : color = 12'he73;
15'b0000101010101101101 : color = 12'he73;
15'b0000101010101101110 : color = 12'he73;
15'b0000101010101101111 : color = 12'he73;
15'b0000101010101110000 : color = 12'he73;
15'b0000101010101110001 : color = 12'he73;
15'b0000101010101110010 : color = 12'he73;
15'b0000101010101110011 : color = 12'he73;
15'b0000101010101110100 : color = 12'he73;
15'b0000101010101110101 : color = 12'he73;
15'b0000101010101110110 : color = 12'he73;
15'b0000101010101110111 : color = 12'he73;
15'b0000101010101111000 : color = 12'he73;
15'b0000101010101111001 : color = 12'he73;
15'b0000101010101111010 : color = 12'he73;
15'b0000101010101111011 : color = 12'he73;
15'b0000101010101111100 : color = 12'he73;
15'b0000101010101111101 : color = 12'he73;
15'b0000101010101111110 : color = 12'he73;
15'b0000101010101111111 : color = 12'he73;
15'b0000101010110000000 : color = 12'he73;
15'b0000101010110000001 : color = 12'he73;
15'b0000101010110000010 : color = 12'he73;
15'b0000101010110000011 : color = 12'he73;
15'b0000101010110000100 : color = 12'he73;
15'b0000101010110000101 : color = 12'he73;
15'b0000101010110000110 : color = 12'he73;
15'b0000101010110000111 : color = 12'he73;
15'b0000101010110001000 : color = 12'he73;
15'b0000101010110001001 : color = 12'he73;
15'b0000101010110001010 : color = 12'he73;
15'b0000101010110001011 : color = 12'he73;
15'b0000101010110001100 : color = 12'he73;
15'b0000101010110001101 : color = 12'he73;
15'b0000101010110001110 : color = 12'he73;
15'b0000101010110001111 : color = 12'he73;
15'b0000101010110010000 : color = 12'he73;
15'b0000101010110010001 : color = 12'he73;
15'b0000101010110010010 : color = 12'he73;
15'b0000101010110010011 : color = 12'he73;
15'b0000101010110010100 : color = 12'he73;
15'b0000101010110010101 : color = 12'he73;
15'b0000101010110010110 : color = 12'he73;
15'b0000101010110010111 : color = 12'he73;
15'b0000101010110011000 : color = 12'he73;
15'b0000101010110011001 : color = 12'he73;
15'b0000101010110011010 : color = 12'he73;
15'b0000101010110011011 : color = 12'he73;
15'b0000101010110011100 : color = 12'he73;
15'b0000101010110011101 : color = 12'he73;
15'b0000101010110011110 : color = 12'he73;
15'b0000101010110011111 : color = 12'he73;
15'b0000101010110100000 : color = 12'he73;
15'b0000101010110100001 : color = 12'he73;
15'b0000101010110100010 : color = 12'he73;
15'b0000101010110100011 : color = 12'he73;
15'b0000101010110100100 : color = 12'he73;
15'b0000101010110100101 : color = 12'he73;
15'b0000101010110100110 : color = 12'he73;
15'b0000101010110100111 : color = 12'he73;
15'b0000101010110101000 : color = 12'he73;
15'b0000101010110101001 : color = 12'he73;
15'b0000101010110101010 : color = 12'he73;
15'b0000101010110101011 : color = 12'he73;
15'b0000101010110101100 : color = 12'he73;
15'b0000101010110101101 : color = 12'he73;
15'b0000101010110101110 : color = 12'he73;
15'b0000101010110101111 : color = 12'he73;
15'b0000101010110110000 : color = 12'he73;
15'b0000101010110110001 : color = 12'he73;
15'b0000101010110110010 : color = 12'he73;
15'b0000101010110110011 : color = 12'he73;
15'b0000101010110110100 : color = 12'he73;
15'b0000101010110110101 : color = 12'he73;
15'b0000101010110110110 : color = 12'he73;
15'b0000101010110110111 : color = 12'he73;
15'b0000101010110111000 : color = 12'he73;
15'b0000101010110111001 : color = 12'he73;
15'b0000101010110111010 : color = 12'he73;
15'b0000101010110111011 : color = 12'he73;
15'b0000101010110111100 : color = 12'he73;
15'b0000101010110111101 : color = 12'he73;
15'b0000101010110111110 : color = 12'he73;
15'b0000101010110111111 : color = 12'he73;
15'b0000101010111000000 : color = 12'he73;
15'b0000101010111000001 : color = 12'he73;
15'b0000101010111000010 : color = 12'he73;
15'b0000101010111000011 : color = 12'he73;
15'b0000101010111000100 : color = 12'he73;
15'b0000101010111000101 : color = 12'he73;
15'b0000101010111000110 : color = 12'he73;
15'b0000101010111000111 : color = 12'he73;
15'b0000101010111001000 : color = 12'he73;
15'b0000101010111001001 : color = 12'he73;
15'b0000101010111001010 : color = 12'he73;
15'b0000101010111001011 : color = 12'he73;
15'b0000101010111001100 : color = 12'he73;
15'b0000101010111001101 : color = 12'he73;
15'b0000101010111001110 : color = 12'he73;
15'b0000101010111001111 : color = 12'he73;
15'b0000101010111010000 : color = 12'he73;
15'b0000101010111010001 : color = 12'he73;
15'b0000101010111010010 : color = 12'he73;
15'b0000101010111010011 : color = 12'he73;
15'b0000101010111010100 : color = 12'he73;
15'b0000101010111010101 : color = 12'he73;
15'b0000101010111010110 : color = 12'he73;
15'b0000101010111010111 : color = 12'he73;
15'b0000101010111011000 : color = 12'he73;
15'b0000101010111011001 : color = 12'he73;
15'b0000101010111011010 : color = 12'he73;
15'b0000101010111011011 : color = 12'he73;
15'b0000101010111011100 : color = 12'he73;
15'b0000101010111011101 : color = 12'he73;
15'b0000101010111011110 : color = 12'he73;
15'b0000101010111011111 : color = 12'he73;
15'b0000101010111100000 : color = 12'he73;
15'b0000101010111100001 : color = 12'he73;
15'b0000101010111100010 : color = 12'he73;
15'b0000101010111100011 : color = 12'he73;
15'b0000101010111100100 : color = 12'he73;
15'b0000101010111100101 : color = 12'he73;
15'b0000101010111100110 : color = 12'he73;
15'b0000101010111100111 : color = 12'he73;
15'b0000101010111101000 : color = 12'he73;
15'b0000101010111101001 : color = 12'he73;
15'b0000101010111101010 : color = 12'he73;
15'b0000101010111101011 : color = 12'he73;
15'b0000101010111101100 : color = 12'he73;
15'b0000101010111101101 : color = 12'he73;
15'b0000101010111101110 : color = 12'he73;
15'b0000101010111101111 : color = 12'he73;
15'b0000101010111110000 : color = 12'he73;
15'b0000101010111110001 : color = 12'he73;
15'b0000101010111110010 : color = 12'he73;
15'b0000101010111110011 : color = 12'he73;
15'b0000101010111110100 : color = 12'he73;
15'b0000101010111110101 : color = 12'he73;
15'b0000101010111110110 : color = 12'he73;
15'b0000101010111110111 : color = 12'he73;
15'b0000101010111111000 : color = 12'he73;
15'b0000101010111111001 : color = 12'he73;
15'b0000101010111111010 : color = 12'he73;
15'b0000101010111111011 : color = 12'he73;
15'b0000101010111111100 : color = 12'he73;
15'b0000101010111111101 : color = 12'he73;
15'b0000101010111111110 : color = 12'he73;
15'b0000101010111111111 : color = 12'he73;
15'b0000101011000000000 : color = 12'he73;
15'b0000101011000000001 : color = 12'he73;
15'b0000101011000000010 : color = 12'he73;
15'b0000101011000000011 : color = 12'he73;
15'b0000101011000000100 : color = 12'he73;
15'b0000101011000000101 : color = 12'he73;
15'b0000101011000000110 : color = 12'he73;
15'b0000101011000000111 : color = 12'he73;
15'b0000101011000001000 : color = 12'he73;
15'b0000101011000001001 : color = 12'he73;
15'b0000101011000001010 : color = 12'he73;
15'b0000101011000001011 : color = 12'he73;
15'b0000101011000001100 : color = 12'he73;
15'b0000101011000001101 : color = 12'he73;
15'b0000101011000001110 : color = 12'he73;
15'b0000101011000001111 : color = 12'he73;
15'b0000101011000010000 : color = 12'he73;
15'b0000101011000010001 : color = 12'he73;
15'b0000101011000010010 : color = 12'he73;
15'b0000101011000010011 : color = 12'he73;
15'b0000101011000010100 : color = 12'he73;
15'b0000101011000010101 : color = 12'he73;
15'b0000101011000010110 : color = 12'he73;
15'b0000101011000010111 : color = 12'he73;
15'b0000101011000011000 : color = 12'he73;
15'b0000101011000011001 : color = 12'he73;
15'b0000101011000011010 : color = 12'he73;
15'b0000101011000011011 : color = 12'he73;
15'b0000101011000011100 : color = 12'he73;
15'b0000101011000011101 : color = 12'he73;
15'b0000101011000011110 : color = 12'he73;
15'b0000101011000011111 : color = 12'he73;
15'b0000101011000100000 : color = 12'he73;
15'b0000101011000100001 : color = 12'he73;
15'b0000101011000100010 : color = 12'he73;
15'b0000101011000100011 : color = 12'he73;
15'b0000101011000100100 : color = 12'he73;
15'b0000101011000100101 : color = 12'he73;
15'b0000101011000100110 : color = 12'he73;
15'b0000101011000100111 : color = 12'he73;
15'b0000101011000101000 : color = 12'he73;
15'b0000101011000101001 : color = 12'he73;
15'b0000101011000101010 : color = 12'he73;
15'b0000101011000101011 : color = 12'he73;
15'b0000101011000101100 : color = 12'he73;
15'b0000101011000101101 : color = 12'he73;
15'b0000101011000101110 : color = 12'he73;
15'b0000101011000101111 : color = 12'he73;
15'b0000101011000110000 : color = 12'he73;
15'b0000101011000110001 : color = 12'he73;
15'b0000101011000110010 : color = 12'he73;
15'b0000101011000110011 : color = 12'he73;
15'b0000101011000110100 : color = 12'he73;
15'b0000101011000110101 : color = 12'he73;
15'b0000101011000110110 : color = 12'he73;
15'b0000101011000110111 : color = 12'he73;
15'b0000101011000111000 : color = 12'he73;
15'b0000101011000111001 : color = 12'he73;
15'b0000101011000111010 : color = 12'he73;
15'b0000101011000111011 : color = 12'he73;
15'b0000101011000111100 : color = 12'he73;
15'b0000101011000111101 : color = 12'he73;
15'b0000101011000111110 : color = 12'he73;
15'b0000101011000111111 : color = 12'he73;
15'b0000101011001000000 : color = 12'he73;
15'b0000101011001000001 : color = 12'he73;
15'b0000101011001000010 : color = 12'he73;
15'b0000101011001000011 : color = 12'he73;
15'b0000101011001000100 : color = 12'he73;
15'b0000101011001000101 : color = 12'he73;
15'b0000101011001000110 : color = 12'he73;
15'b0000101011001000111 : color = 12'he73;
15'b0000101011001001000 : color = 12'he73;
15'b0000101011001001001 : color = 12'he73;
15'b0000101011001001010 : color = 12'he73;
15'b0000101011001001011 : color = 12'he73;
15'b0000101011001001100 : color = 12'he73;
15'b0000101011001001101 : color = 12'he73;
15'b0000101011001001110 : color = 12'he73;
15'b0000101011001001111 : color = 12'he73;
15'b0000101011001010000 : color = 12'he73;
15'b0000101011001010001 : color = 12'he73;
15'b0000101011001010010 : color = 12'he73;
15'b0000101011001010011 : color = 12'he73;
15'b0000101011001010100 : color = 12'he73;
15'b0000101011001010101 : color = 12'he73;
15'b0000101011001010110 : color = 12'he73;
15'b0000101011001010111 : color = 12'he73;
15'b0000101011001011000 : color = 12'he73;
15'b0000101011001011001 : color = 12'he73;
15'b0000101011001011010 : color = 12'he73;
15'b0000101011001011011 : color = 12'he73;
15'b0000101011001011100 : color = 12'he73;
15'b0000101011001011101 : color = 12'he73;
15'b0000101011001011110 : color = 12'he73;
15'b0000101011001011111 : color = 12'he73;
15'b0000101011001100000 : color = 12'he73;
15'b0000101011001100001 : color = 12'he73;
15'b0000101011001100010 : color = 12'he73;
15'b0000101011001100011 : color = 12'he73;
15'b0000101011001100100 : color = 12'he73;
15'b0000101011001100101 : color = 12'he73;
15'b0000101011001100110 : color = 12'he73;
15'b0000101011001100111 : color = 12'he73;
15'b0000101011001101000 : color = 12'he73;
15'b0000101011001101001 : color = 12'he73;
15'b0000101011001101010 : color = 12'he73;
15'b0000101011001101011 : color = 12'he73;
15'b0000101011001101100 : color = 12'he73;
15'b0000101011001101101 : color = 12'he73;
15'b0000101011001101110 : color = 12'he73;
15'b0000101011001101111 : color = 12'he73;
15'b0000101011001110000 : color = 12'he73;
15'b0000101011001110001 : color = 12'he73;
15'b0000101011001110010 : color = 12'he73;
15'b0000101011001110011 : color = 12'he73;
15'b0000101011001110100 : color = 12'he73;
15'b0000101011001110101 : color = 12'he73;
15'b0000101011001110110 : color = 12'he73;
15'b0000101011001110111 : color = 12'he73;
15'b0000101011001111000 : color = 12'he73;
15'b0000101011001111001 : color = 12'he73;
15'b0000101011001111010 : color = 12'he73;
15'b0000101011001111011 : color = 12'he73;
15'b0000101011001111100 : color = 12'he73;
15'b0000101011001111101 : color = 12'he73;
15'b0000101011001111110 : color = 12'he73;
15'b0000101011001111111 : color = 12'he73;
15'b0000101011010000000 : color = 12'he73;
15'b0000101011010000001 : color = 12'he73;
15'b0000101011010000010 : color = 12'he73;
15'b0000101011010000011 : color = 12'he73;
15'b0000101011010000100 : color = 12'he73;
15'b0000101011010000101 : color = 12'he73;
15'b0000101011010000110 : color = 12'he73;
15'b0000101011010000111 : color = 12'he73;
15'b0000101011010001000 : color = 12'he73;
15'b0000101011010001001 : color = 12'he73;
15'b0000101011010001010 : color = 12'he73;
15'b0000101011010001011 : color = 12'he73;
15'b0000101011010001100 : color = 12'he73;
15'b0000101011010001101 : color = 12'he73;
15'b0000101011010001110 : color = 12'he73;
15'b0000101011010001111 : color = 12'he73;
15'b0000101011010010000 : color = 12'he73;
15'b0000101011010010001 : color = 12'he73;
15'b0000101011010010010 : color = 12'he73;
15'b0000101011010010011 : color = 12'he73;
15'b0000101011010010100 : color = 12'he73;
15'b0000101011010010101 : color = 12'he73;
15'b0000101011010010110 : color = 12'he73;
15'b0000101011010010111 : color = 12'he73;
15'b0000101011010011000 : color = 12'he73;
15'b0000101011010011001 : color = 12'he73;
15'b0000101011010011010 : color = 12'he73;
15'b0000101011010011011 : color = 12'he73;
15'b0000101011010011100 : color = 12'he73;
15'b0000101011010011101 : color = 12'he73;
15'b0000101011010011110 : color = 12'he73;
15'b0000101011010011111 : color = 12'he73;
15'b0000101011010100000 : color = 12'he73;
15'b0000101011010100001 : color = 12'he73;
15'b0000101011010100010 : color = 12'he73;
15'b0000101011010100011 : color = 12'he73;
15'b0000101010011100010 : color = 12'he73;
15'b0000101010011100011 : color = 12'he73;
15'b0000101010011100100 : color = 12'he73;
15'b0000101010011100101 : color = 12'he73;
15'b0000101010011100110 : color = 12'he73;
15'b0000101010011100111 : color = 12'he73;
15'b0000101010011101000 : color = 12'he73;
15'b0000101010011101001 : color = 12'he73;
15'b0000101010011101010 : color = 12'he73;
15'b0000101010011101011 : color = 12'he73;
15'b0000101010011101100 : color = 12'he73;
15'b0000101010011101101 : color = 12'he73;
15'b0000101010011101110 : color = 12'he73;
15'b0000101010011101111 : color = 12'he73;
15'b0000101010011110000 : color = 12'he73;
15'b0000101010011110001 : color = 12'he73;
15'b0000101010011110010 : color = 12'he73;
15'b0000101010011110011 : color = 12'he73;
15'b0000101010011110100 : color = 12'he73;
15'b0000101010011110101 : color = 12'he73;
15'b0000101010011110110 : color = 12'he73;
15'b0000101010011110111 : color = 12'he73;
15'b0000101010011111000 : color = 12'he73;
15'b0000101010011111001 : color = 12'he73;
15'b0000101010011111010 : color = 12'he73;
15'b0000101010011111011 : color = 12'he73;
15'b0000101010011111100 : color = 12'he73;
15'b0000101010011111101 : color = 12'he73;
15'b0000101010011111110 : color = 12'he73;
15'b0000101010011111111 : color = 12'he73;
15'b0000101010100000000 : color = 12'he73;
15'b0000101010100000001 : color = 12'he73;
15'b0000101010100000010 : color = 12'he73;
15'b0000101010100000011 : color = 12'he73;
15'b0000101010100000100 : color = 12'he73;
15'b0000101010100000101 : color = 12'he73;
15'b0000101010100000110 : color = 12'he73;
15'b0000101010100000111 : color = 12'he73;
15'b0000101010100001000 : color = 12'he73;
15'b0000101010100001001 : color = 12'he73;
15'b0000101010100001010 : color = 12'he73;
15'b0000101010100001011 : color = 12'he73;
15'b0000101010100001100 : color = 12'he73;
15'b0000101010100001101 : color = 12'he73;
15'b0000101010100001110 : color = 12'he73;
15'b0000101010100001111 : color = 12'he73;
15'b0000101010100010000 : color = 12'he73;
15'b0000101010100010001 : color = 12'he73;
15'b0000101010100010010 : color = 12'he73;
15'b0000101010100010011 : color = 12'he73;
15'b0000101010100010100 : color = 12'he73;
15'b0000101010100010101 : color = 12'he73;
15'b0000101010100010110 : color = 12'he73;
15'b0000101010100010111 : color = 12'he73;
15'b0000101010100011000 : color = 12'he73;
15'b0000101010100011001 : color = 12'he73;
15'b0000101010100011010 : color = 12'he73;
15'b0000101010100011011 : color = 12'he73;
15'b0000101010100011100 : color = 12'he73;
15'b0000101010100011101 : color = 12'he73;
15'b0000101010100011110 : color = 12'he73;
15'b0000101010100011111 : color = 12'he73;
15'b0000101010100100000 : color = 12'he73;
15'b0000101010100100001 : color = 12'he73;
15'b0000101010100100010 : color = 12'he73;
15'b0000101010100100011 : color = 12'he73;
15'b0000101010100100100 : color = 12'he73;
15'b0000101010100100101 : color = 12'he73;
15'b0000101010100100110 : color = 12'he73;
15'b0000101010100100111 : color = 12'he73;
15'b0000101010100101000 : color = 12'he73;
15'b0000101010100101001 : color = 12'he73;
15'b0000101010100101010 : color = 12'he73;
15'b0000101010100101011 : color = 12'he73;
15'b0000101010100101100 : color = 12'he73;
15'b0000101010100101101 : color = 12'he73;
15'b0000101010100101110 : color = 12'he73;
15'b0000101010100101111 : color = 12'he73;
15'b0000101010100110000 : color = 12'he73;
15'b0000101010100110001 : color = 12'he73;
15'b0000101010100110010 : color = 12'he73;
15'b0000101010100110011 : color = 12'he73;
15'b0000101010100110100 : color = 12'he73;
15'b0000101010100110101 : color = 12'he73;
15'b0000101010100110110 : color = 12'he73;
15'b0000101010100110111 : color = 12'he73;
15'b0000101010100111000 : color = 12'he73;
15'b0000101010100111001 : color = 12'he73;
15'b0000101010100111010 : color = 12'he73;
15'b0000101010100111011 : color = 12'he73;
15'b0000101010100111100 : color = 12'he73;
15'b0000101010100111101 : color = 12'he73;
15'b0000101010100111110 : color = 12'he73;
15'b0000101010100111111 : color = 12'he73;
15'b0000101010101000000 : color = 12'he73;
15'b0000101010101000001 : color = 12'he73;
15'b0000101010101000010 : color = 12'he73;
15'b0000101010101000011 : color = 12'he73;
15'b0000101010101000100 : color = 12'he73;
15'b0000101010101000101 : color = 12'he73;
15'b0000101010101000110 : color = 12'he73;
15'b0000101010101000111 : color = 12'he73;
15'b0000101010101001000 : color = 12'he73;
15'b0000101010101001001 : color = 12'he73;
15'b0000101010101001010 : color = 12'he73;
15'b0000101010101001011 : color = 12'he73;
15'b0000101010101001100 : color = 12'he73;
15'b0000101010101001101 : color = 12'he73;
15'b0000101010101001110 : color = 12'he73;
15'b0000101010101001111 : color = 12'he73;
15'b0000101010101010000 : color = 12'he73;
15'b0000101010101010001 : color = 12'he73;
15'b0000101010101010010 : color = 12'he73;
15'b0000101010101010011 : color = 12'he73;
15'b0000101010101010100 : color = 12'he73;
15'b0000101010101010101 : color = 12'he73;
15'b0000101010101010110 : color = 12'he73;
15'b0000101010101010111 : color = 12'he73;
15'b0000101010101011000 : color = 12'he73;
15'b0000101010101011001 : color = 12'he73;
15'b0000101010101011010 : color = 12'he73;
15'b0000101010101011011 : color = 12'he73;
15'b0000101010101011100 : color = 12'he73;
15'b0000101010101011101 : color = 12'he73;
15'b0000101010101011110 : color = 12'he73;
15'b0000101010101011111 : color = 12'he73;
15'b0000101010101100000 : color = 12'he73;
15'b0000101010101100001 : color = 12'he73;
15'b0000101010101100010 : color = 12'he73;
15'b0000101010101100011 : color = 12'he73;
15'b0000101010101100100 : color = 12'he73;
15'b0000101010101100101 : color = 12'he73;
15'b0000101010101100110 : color = 12'he73;
15'b0000101010101100111 : color = 12'he73;
15'b0000101010101101000 : color = 12'he73;
15'b0000101010101101001 : color = 12'he73;
15'b0000101010101101010 : color = 12'he73;
15'b0000101010101101011 : color = 12'he73;
15'b0000101010101101100 : color = 12'he73;
15'b0000101010101101101 : color = 12'he73;
15'b0000101010101101110 : color = 12'he73;
15'b0000101010101101111 : color = 12'he73;
15'b0000101010101110000 : color = 12'he73;
15'b0000101010101110001 : color = 12'he73;
15'b0000101010101110010 : color = 12'he73;
15'b0000101010101110011 : color = 12'he73;
15'b0000101010101110100 : color = 12'he73;
15'b0000101010101110101 : color = 12'he73;
15'b0000101010101110110 : color = 12'he73;
15'b0000101010101110111 : color = 12'he73;
15'b0000101010101111000 : color = 12'he73;
15'b0000101010101111001 : color = 12'he73;
15'b0000101010101111010 : color = 12'he73;
15'b0000101010101111011 : color = 12'he73;
15'b0000101010101111100 : color = 12'he73;
15'b0000101010101111101 : color = 12'he73;
15'b0000101010101111110 : color = 12'he73;
15'b0000101010101111111 : color = 12'he73;
15'b0000101010110000000 : color = 12'he73;
15'b0000101010110000001 : color = 12'he73;
15'b0000101010110000010 : color = 12'he73;
15'b0000101010110000011 : color = 12'he73;
15'b0000101010110000100 : color = 12'he73;
15'b0000101010110000101 : color = 12'he73;
15'b0000101010110000110 : color = 12'he73;
15'b0000101010110000111 : color = 12'he73;
15'b0000101010110001000 : color = 12'he73;
15'b0000101010110001001 : color = 12'he73;
15'b0000101010110001010 : color = 12'he73;
15'b0000101010110001011 : color = 12'he73;
15'b0000101010110001100 : color = 12'he73;
15'b0000101010110001101 : color = 12'he73;
15'b0000101010110001110 : color = 12'he73;
15'b0000101010110001111 : color = 12'he73;
15'b0000101010110010000 : color = 12'he73;
15'b0000101010110010001 : color = 12'he73;
15'b0000101010110010010 : color = 12'he73;
15'b0000101010110010011 : color = 12'he73;
15'b0000101010110010100 : color = 12'he73;
15'b0000101010110010101 : color = 12'he73;
15'b0000101010110010110 : color = 12'he73;
15'b0000101010110010111 : color = 12'he73;
15'b0000101010110011000 : color = 12'he73;
15'b0000101010110011001 : color = 12'he73;
15'b0000101010110011010 : color = 12'he73;
15'b0000101010110011011 : color = 12'he73;
15'b0000101010110011100 : color = 12'he73;
15'b0000101010110011101 : color = 12'he73;
15'b0000101010110011110 : color = 12'he73;
15'b0000101010110011111 : color = 12'he73;
15'b0000101010110100000 : color = 12'he73;
15'b0000101010110100001 : color = 12'he73;
15'b0000101010110100010 : color = 12'he73;
15'b0000101010110100011 : color = 12'he73;
15'b0000101010110100100 : color = 12'he73;
15'b0000101010110100101 : color = 12'he73;
15'b0000101010110100110 : color = 12'he73;
15'b0000101010110100111 : color = 12'he73;
15'b0000101010110101000 : color = 12'he73;
15'b0000101010110101001 : color = 12'he73;
15'b0000101010110101010 : color = 12'he73;
15'b0000101010110101011 : color = 12'he73;
15'b0000101010110101100 : color = 12'he73;
15'b0000101010110101101 : color = 12'he73;
15'b0000101010110101110 : color = 12'he73;
15'b0000101010110101111 : color = 12'he73;
15'b0000101010110110000 : color = 12'he73;
15'b0000101010110110001 : color = 12'he73;
15'b0000101010110110010 : color = 12'he73;
15'b0000101010110110011 : color = 12'he73;
15'b0000101010110110100 : color = 12'he73;
15'b0000101010110110101 : color = 12'he73;
15'b0000101010110110110 : color = 12'he73;
15'b0000101010110110111 : color = 12'he73;
15'b0000101010110111000 : color = 12'he73;
15'b0000101010110111001 : color = 12'he73;
15'b0000101010110111010 : color = 12'he73;
15'b0000101010110111011 : color = 12'he73;
15'b0000101010110111100 : color = 12'he73;
15'b0000101010110111101 : color = 12'he73;
15'b0000101010110111110 : color = 12'he73;
15'b0000101010110111111 : color = 12'he73;
15'b0000101010111000000 : color = 12'he73;
15'b0000101010111000001 : color = 12'he73;
15'b0000101010111000010 : color = 12'he73;
15'b0000101010111000011 : color = 12'he73;
15'b0000101010111000100 : color = 12'he73;
15'b0000101010111000101 : color = 12'he73;
15'b0000101010111000110 : color = 12'he73;
15'b0000101010111000111 : color = 12'he73;
15'b0000101010111001000 : color = 12'he73;
15'b0000101010111001001 : color = 12'he73;
15'b0000101010111001010 : color = 12'he73;
15'b0000101010111001011 : color = 12'he73;
15'b0000101010111001100 : color = 12'he73;
15'b0000101010111001101 : color = 12'he73;
15'b0000101010111001110 : color = 12'he73;
15'b0000101010111001111 : color = 12'he73;
15'b0000101010111010000 : color = 12'he73;
15'b0000101010111010001 : color = 12'he73;
15'b0000101010111010010 : color = 12'he73;
15'b0000101010111010011 : color = 12'he73;
15'b0000101010111010100 : color = 12'he73;
15'b0000101010111010101 : color = 12'he73;
15'b0000101010111010110 : color = 12'he73;
15'b0000101010111010111 : color = 12'he73;
15'b0000101010111011000 : color = 12'he73;
15'b0000101010111011001 : color = 12'he73;
15'b0000101010111011010 : color = 12'he73;
15'b0000101010111011011 : color = 12'he73;
15'b0000101010111011100 : color = 12'he73;
15'b0000101010111011101 : color = 12'he73;
15'b0000101010111011110 : color = 12'he73;
15'b0000101010111011111 : color = 12'he73;
15'b0000101010111100000 : color = 12'he73;
15'b0000101010111100001 : color = 12'he73;
15'b0000101010111100010 : color = 12'he73;
15'b0000101010111100011 : color = 12'he73;
15'b0000101010111100100 : color = 12'he73;
15'b0000101010111100101 : color = 12'he73;
15'b0000101010111100110 : color = 12'he73;
15'b0000101010111100111 : color = 12'he73;
15'b0000101010111101000 : color = 12'he73;
15'b0000101010111101001 : color = 12'he73;
15'b0000101010111101010 : color = 12'he73;
15'b0000101010111101011 : color = 12'he73;
15'b0000101010111101100 : color = 12'he73;
15'b0000101010111101101 : color = 12'he73;
15'b0000101010111101110 : color = 12'he73;
15'b0000101010111101111 : color = 12'he73;
15'b0000101010111110000 : color = 12'he73;
15'b0000101010111110001 : color = 12'he73;
15'b0000101010111110010 : color = 12'he73;
15'b0000101010111110011 : color = 12'he73;
15'b0000101010111110100 : color = 12'he73;
15'b0000101010111110101 : color = 12'he73;
15'b0000101010111110110 : color = 12'he73;
15'b0000101010111110111 : color = 12'he73;
15'b0000101010111111000 : color = 12'he73;
15'b0000101010111111001 : color = 12'he73;
15'b0000101010111111010 : color = 12'he73;
15'b0000101010111111011 : color = 12'he73;
15'b0000101010111111100 : color = 12'he73;
15'b0000101010111111101 : color = 12'he73;
15'b0000101010111111110 : color = 12'he73;
15'b0000101010111111111 : color = 12'he73;
15'b0000101011000000000 : color = 12'he73;
15'b0000101011000000001 : color = 12'he73;
15'b0000101011000000010 : color = 12'he73;
15'b0000101011000000011 : color = 12'he73;
15'b0000101011000000100 : color = 12'he73;
15'b0000101011000000101 : color = 12'he73;
15'b0000101011000000110 : color = 12'he73;
15'b0000101011000000111 : color = 12'he73;
15'b0000101011000001000 : color = 12'he73;
15'b0000101011000001001 : color = 12'he73;
15'b0000101011000001010 : color = 12'he73;
15'b0000101011000001011 : color = 12'he73;
15'b0000101011000001100 : color = 12'he73;
15'b0000101011000001101 : color = 12'he73;
15'b0000101011000001110 : color = 12'he73;
15'b0000101011000001111 : color = 12'he73;
15'b0000101011000010000 : color = 12'he73;
15'b0000101011000010001 : color = 12'he73;
15'b0000101011000010010 : color = 12'he73;
15'b0000101011000010011 : color = 12'he73;
15'b0000101011000010100 : color = 12'he73;
15'b0000101011000010101 : color = 12'he73;
15'b0000101011000010110 : color = 12'he73;
15'b0000101011000010111 : color = 12'he73;
15'b0000101011000011000 : color = 12'he73;
15'b0000101011000011001 : color = 12'he73;
15'b0000101011000011010 : color = 12'he73;
15'b0000101011000011011 : color = 12'he73;
15'b0000101011000011100 : color = 12'he73;
15'b0000101011000011101 : color = 12'he73;
15'b0000101011000011110 : color = 12'he73;
15'b0000101011000011111 : color = 12'he73;
15'b0000101011000100000 : color = 12'he73;
15'b0000101011000100001 : color = 12'he73;
15'b0000101011000100010 : color = 12'he73;
15'b0000101011000100011 : color = 12'he73;
15'b0000101011000100100 : color = 12'he73;
15'b0000101011000100101 : color = 12'he73;
15'b0000101011000100110 : color = 12'he73;
15'b0000101011000100111 : color = 12'he73;
15'b0000101011000101000 : color = 12'he73;
15'b0000101011000101001 : color = 12'he73;
15'b0000101011000101010 : color = 12'he73;
15'b0000101011000101011 : color = 12'he73;
15'b0000101011000101100 : color = 12'he73;
15'b0000101011000101101 : color = 12'he73;
15'b0000101011000101110 : color = 12'he73;
15'b0000101011000101111 : color = 12'he73;
15'b0000101011000110000 : color = 12'he73;
15'b0000101011000110001 : color = 12'he73;
15'b0000101011000110010 : color = 12'he73;
15'b0000101011000110011 : color = 12'he73;
15'b0000101011000110100 : color = 12'he73;
15'b0000101011000110101 : color = 12'he73;
15'b0000101011000110110 : color = 12'he73;
15'b0000101011000110111 : color = 12'he73;
15'b0000101011000111000 : color = 12'he73;
15'b0000101011000111001 : color = 12'he73;
15'b0000101011000111010 : color = 12'he73;
15'b0000101011000111011 : color = 12'he73;
15'b0000101011000111100 : color = 12'he73;
15'b0000101011000111101 : color = 12'he73;
15'b0000101011000111110 : color = 12'he73;
15'b0000101011000111111 : color = 12'he73;
15'b0000101011001000000 : color = 12'he73;
15'b0000101011001000001 : color = 12'he73;
15'b0000101011001000010 : color = 12'he73;
15'b0000101011001000011 : color = 12'he73;
15'b0000101011001000100 : color = 12'he73;
15'b0000101011001000101 : color = 12'he73;
15'b0000101011001000110 : color = 12'he73;
15'b0000101011001000111 : color = 12'he73;
15'b0000101011001001000 : color = 12'he73;
15'b0000101011001001001 : color = 12'he73;
15'b0000101011001001010 : color = 12'he73;
15'b0000101011001001011 : color = 12'he73;
15'b0000101011001001100 : color = 12'he73;
15'b0000101011001001101 : color = 12'he73;
15'b0000101011001001110 : color = 12'he73;
15'b0000101011001001111 : color = 12'he73;
15'b0000101011001010000 : color = 12'he73;
15'b0000101011001010001 : color = 12'he73;
15'b0000101011001010010 : color = 12'he73;
15'b0000101011001010011 : color = 12'he73;
15'b0000101011001010100 : color = 12'he73;
15'b0000101011001010101 : color = 12'he73;
15'b0000101011001010110 : color = 12'he73;
15'b0000101011001010111 : color = 12'he73;
15'b0000101011001011000 : color = 12'he73;
15'b0000101011001011001 : color = 12'he73;
15'b0000101011001011010 : color = 12'he73;
15'b0000101011001011011 : color = 12'he73;
15'b0000101011001011100 : color = 12'he73;
15'b0000101011001011101 : color = 12'he73;
15'b0000101011001011110 : color = 12'he73;
15'b0000101011001011111 : color = 12'he73;
15'b0000101011001100000 : color = 12'he73;
15'b0000101011001100001 : color = 12'he73;
15'b0000101011001100010 : color = 12'he73;
15'b0000101011001100011 : color = 12'he73;
15'b0000101011001100100 : color = 12'he73;
15'b0000101011001100101 : color = 12'he73;
15'b0000101011001100110 : color = 12'he73;
15'b0000101011001100111 : color = 12'he73;
15'b0000101011001101000 : color = 12'he73;
15'b0000101011001101001 : color = 12'he73;
15'b0000101011001101010 : color = 12'he73;
15'b0000101011001101011 : color = 12'he73;
15'b0000101011001101100 : color = 12'he73;
15'b0000101011001101101 : color = 12'he73;
15'b0000101011001101110 : color = 12'he73;
15'b0000101011001101111 : color = 12'he73;
15'b0000101011001110000 : color = 12'he73;
15'b0000101011001110001 : color = 12'he73;
15'b0000101011001110010 : color = 12'he73;
15'b0000101011001110011 : color = 12'he73;
15'b0000101011001110100 : color = 12'he73;
15'b0000101011001110101 : color = 12'he73;
15'b0000101011001110110 : color = 12'he73;
15'b0000101011001110111 : color = 12'he73;
15'b0000101011001111000 : color = 12'he73;
15'b0000101011001111001 : color = 12'he73;
15'b0000101011001111010 : color = 12'he73;
15'b0000101011001111011 : color = 12'he73;
15'b0000101011001111100 : color = 12'he73;
15'b0000101011001111101 : color = 12'he73;
15'b0000101011001111110 : color = 12'he73;
15'b0000101011001111111 : color = 12'he73;
15'b0000101011010000000 : color = 12'he73;
15'b0000101011010000001 : color = 12'he73;
15'b0000101011010000010 : color = 12'he73;
15'b0000101011010000011 : color = 12'he73;
15'b0000101011010000100 : color = 12'he73;
15'b0000101011010000101 : color = 12'he73;
15'b0000101011010000110 : color = 12'he73;
15'b0000101011010000111 : color = 12'he73;
15'b0000101011010001000 : color = 12'he73;
15'b0000101011010001001 : color = 12'he73;
15'b0000101011010001010 : color = 12'he73;
15'b0000101011010001011 : color = 12'he73;
15'b0000101011010001100 : color = 12'he73;
15'b0000101011010001101 : color = 12'he73;
15'b0000101011010001110 : color = 12'he73;
15'b0000101011010001111 : color = 12'he73;
15'b0000101011010010000 : color = 12'he73;
15'b0000101011010010001 : color = 12'he73;
15'b0000101011010010010 : color = 12'he73;
15'b0000101011010010011 : color = 12'he73;
15'b0000101011010010100 : color = 12'he73;
15'b0000101011010010101 : color = 12'he73;
15'b0000101011010010110 : color = 12'he73;
15'b0000101011010010111 : color = 12'he73;
15'b0000101011010011000 : color = 12'he73;
15'b0000101011010011001 : color = 12'he73;
15'b0000101011010011010 : color = 12'he73;
15'b0000101011010011011 : color = 12'he73;
15'b0000101011010011100 : color = 12'he73;
15'b0000101011010011101 : color = 12'he73;
15'b0000101011010011110 : color = 12'he73;
15'b0000101011010011111 : color = 12'he73;
15'b0000101011010100000 : color = 12'he73;
15'b0000101011010100001 : color = 12'he73;
15'b0000101011010100010 : color = 12'he73;
15'b0000101011010100011 : color = 12'he73;
15'b0000101011010100100 : color = 12'he73;
15'b0000101011010100101 : color = 12'he73;
15'b0000101011010100110 : color = 12'he73;
15'b0000101011010100111 : color = 12'he73;
15'b0000101011010101000 : color = 12'he73;
15'b0000101011010101001 : color = 12'he73;
15'b0000101011010101010 : color = 12'he73;
15'b0000101011010101011 : color = 12'he73;
15'b0000101011010101100 : color = 12'he73;
15'b0000101011010101101 : color = 12'he73;
15'b0000101011010101110 : color = 12'he73;
15'b0000101011010101111 : color = 12'he73;
15'b0000101011010110000 : color = 12'he73;
15'b0000101011010110001 : color = 12'he73;
15'b0000101011010110010 : color = 12'he73;
15'b0000101011010110011 : color = 12'he73;
15'b0000101011010110100 : color = 12'he73;
15'b0000101011010110101 : color = 12'he73;
15'b0000101011010110110 : color = 12'he73;
15'b0000101011010110111 : color = 12'he73;
15'b0000101011010111000 : color = 12'he73;
15'b0000101011010111001 : color = 12'he73;
15'b0000101011010111010 : color = 12'he73;
15'b0000101011010111011 : color = 12'he73;
15'b0000101011010111100 : color = 12'he73;
15'b0000101011010111101 : color = 12'he73;
15'b0000101011010111110 : color = 12'he73;
15'b0000101011010111111 : color = 12'he73;
15'b0000101011011000000 : color = 12'he73;
15'b0000101011011000001 : color = 12'he73;
15'b0000101011011000010 : color = 12'he73;
15'b0000101011011000011 : color = 12'he73;
15'b0000101011011000100 : color = 12'he73;
15'b0000101011011000101 : color = 12'he73;
15'b0000101011011000110 : color = 12'he73;
15'b0000101011011000111 : color = 12'he73;
15'b0000101011011001000 : color = 12'he73;
15'b0000101011011001001 : color = 12'he73;
15'b0000101011011001010 : color = 12'he73;
15'b0000101011011001011 : color = 12'he73;
15'b0000101011011001100 : color = 12'he73;

default : color = 12'hzzz;
endcase
end
end
endmodule
